module top (
        input wire        sys_clk,
        input wire        sys_rst_n,
        input wire        sink_star,
        input wire        sink_stop,
        input wire [3:0] sink,

    output wire [ 4:0] iter,
    output wire [63:0] data_decode,
        output wire        data_en,
        output wire        buffer_full


    );

    // buffer模块
    wire [3:0] rr_data       [532:0];
    wire [6:0] buffer_addr;  // ram_llr 内部索引地址
    wire [1:0] flag_buffer_in;
    wire        buffer_wr_en;
    wire        flag_org_write_end;

    // 控制模块
    wire        flag_first_store;
    wire        flag_org_read_start;
    wire [23:0] flag_org_read_end;
    wire        flag_CFU_start;
    wire [3:0] flag_CFU_end;
    wire        flag_VFU_start;
    wire [23:0] flag_VFU_end;
    wire        flag_judge_start;
    wire        flag_judge_end;
    wire        flag_org_update;
    wire        flag_serial;

    // 误差错误统计
    wire [ 6:0] H_sum;

    // combine_ram_llr模块
    wire [ 7:0] org_addr     [532:0];  // 533路 llr 数据对应的地址信息，每一路有 7 位的地址
    wire [532:0] org_wr_en;
    wire [2:0] org_data     [532:0];  //有533路原始数据输出到H存储ram中

    // 判决接收
    wire [63:0] bit_data     [532:0];



    // CFU，VFU，ram 之间的连接线
    `include "CV_pin_H_QC_N68224_K65536_R0.96_z128.txt"
    /* wire	[15:0]	ram_CFU_data_1_2;
    wire	[15:0]	CFU_data_1_2;
    wire	[15:0]	ram_VFU_data_1_2;
    wire	[15:0]	VFU_data_1_2;

    wire	[4:0]	CFU_addr_1;//12路
    wire			CFU_wr_en_1;
    wire			CFU_re_en_1;

    wire	[4:0]	VFU_addr_1;//24路
    wire			VFU_wr_en_1;
    wire			VFU_re_en_1; */


    buffer_in #(
                  .QNT_BIT           (3),
                  .QC_LDPC_COL_COUNT (533),
                  .QC_LDPC_BLOCK_SIZE(64)
              ) u_buffer_in (
                  .sys_clk          (sys_clk),
                  .sys_rst_n        (sys_rst_n),
                  .sink_star        (sink_star),
                  .sink_stop        (sink_stop),
                  .sink             (sink),
                  .flag_org_update  (flag_org_update),

                  .buffer_wr_en  (buffer_wr_en),

                   .rr_data_1  (rr_data[0 ]),
                   .rr_data_2  (rr_data[1 ]),
                   .rr_data_3  (rr_data[2 ]),
                   .rr_data_4  (rr_data[3 ]),
                   .rr_data_5  (rr_data[4 ]),
                   .rr_data_6  (rr_data[5 ]),
                   .rr_data_7  (rr_data[6 ]),
                   .rr_data_8  (rr_data[7 ]),
                   .rr_data_9  (rr_data[8 ]),
                   .rr_data_10 (rr_data[9 ]),
                   .rr_data_11 (rr_data[10]),
                   .rr_data_12 (rr_data[11]),
                   .rr_data_13 (rr_data[12]),
                   .rr_data_14 (rr_data[13]),
                   .rr_data_15 (rr_data[14]),
                   .rr_data_16 (rr_data[15]),
                   .rr_data_17 (rr_data[16]),
                   .rr_data_18 (rr_data[17]),
                   .rr_data_19 (rr_data[18]),
                   .rr_data_20 (rr_data[19]),
                   .rr_data_21 (rr_data[20]),
                   .rr_data_22 (rr_data[21]),
                   .rr_data_23 (rr_data[22]),
                   .rr_data_24 (rr_data[23]),
                   .rr_data_25 (rr_data[24]),
                   .rr_data_26 (rr_data[25]),
                   .rr_data_27 (rr_data[26]),
                   .rr_data_28 (rr_data[27]),
                   .rr_data_29 (rr_data[28]),
                   .rr_data_30 (rr_data[29]),
                   .rr_data_31 (rr_data[30]),
                   .rr_data_32 (rr_data[31]),
                   .rr_data_33 (rr_data[32]),
                   .rr_data_34 (rr_data[33]),
                   .rr_data_35 (rr_data[34]),
                   .rr_data_36 (rr_data[35]),
                   .rr_data_37 (rr_data[36]),
                   .rr_data_38 (rr_data[37]),
                   .rr_data_39 (rr_data[38]),
                   .rr_data_40 (rr_data[39]),
                   .rr_data_41 (rr_data[40]),
                   .rr_data_42 (rr_data[41]),
                   .rr_data_43 (rr_data[42]),
                   .rr_data_44 (rr_data[43]),
                   .rr_data_45 (rr_data[44]),
                   .rr_data_46 (rr_data[45]),
                   .rr_data_47 (rr_data[46]),
                   .rr_data_48 (rr_data[47]),
                   .rr_data_49 (rr_data[48]),
                   .rr_data_50 (rr_data[49]),
                   .rr_data_51 (rr_data[50]),
                   .rr_data_52 (rr_data[51]),
                   .rr_data_53 (rr_data[52]),
                   .rr_data_54 (rr_data[53]),
                   .rr_data_55 (rr_data[54]),
                   .rr_data_56 (rr_data[55]),
                   .rr_data_57 (rr_data[56]),
                   .rr_data_58 (rr_data[57]),
                   .rr_data_59 (rr_data[58]),
                   .rr_data_60 (rr_data[59]),
                   .rr_data_61 (rr_data[60]),
                   .rr_data_62 (rr_data[61]),
                   .rr_data_63 (rr_data[62]),
                   .rr_data_64 (rr_data[63]),
                   .rr_data_65 (rr_data[64]),
                   .rr_data_66 (rr_data[65]),
                   .rr_data_67 (rr_data[66]),
                   .rr_data_68 (rr_data[67]),
                   .rr_data_69 (rr_data[68]),
                   .rr_data_70 (rr_data[69]),
                   .rr_data_71 (rr_data[70]),
                   .rr_data_72 (rr_data[71]),
                   .rr_data_73 (rr_data[72]),
                   .rr_data_74 (rr_data[73]),
                   .rr_data_75 (rr_data[74]),
                   .rr_data_76 (rr_data[75]),
                   .rr_data_77 (rr_data[76]),
                   .rr_data_78 (rr_data[77]),
                   .rr_data_79 (rr_data[78]),
                   .rr_data_80 (rr_data[79]),
                   .rr_data_81 (rr_data[80]),
                   .rr_data_82 (rr_data[81]),
                   .rr_data_83 (rr_data[82]),
                   .rr_data_84 (rr_data[83]),
                   .rr_data_85 (rr_data[84]),
                   .rr_data_86 (rr_data[85]),
                   .rr_data_87 (rr_data[86]),
                   .rr_data_88 (rr_data[87]),
                   .rr_data_89 (rr_data[88]),
                   .rr_data_90 (rr_data[89]),
                   .rr_data_91 (rr_data[90]),
                   .rr_data_92 (rr_data[91]),
                   .rr_data_93 (rr_data[92]),
                   .rr_data_94 (rr_data[93]),
                   .rr_data_95 (rr_data[94]),
                   .rr_data_96 (rr_data[95]),
                   .rr_data_97 (rr_data[96]),
                   .rr_data_98 (rr_data[97]),
                   .rr_data_99 (rr_data[98]),
                   .rr_data_100(rr_data[99]),
                   .rr_data_101(rr_data[100]),
                   .rr_data_102(rr_data[101]),
                   .rr_data_103(rr_data[102]),
                   .rr_data_104(rr_data[103]),
                   .rr_data_105(rr_data[104]),
                   .rr_data_106(rr_data[105]),
                   .rr_data_107(rr_data[106]),
                   .rr_data_108(rr_data[107]),
                   .rr_data_109(rr_data[108]),
                   .rr_data_110(rr_data[109]),
                   .rr_data_111(rr_data[110]),
                   .rr_data_112(rr_data[111]),
                   .rr_data_113(rr_data[112]),
                   .rr_data_114(rr_data[113]),
                   .rr_data_115(rr_data[114]),
                   .rr_data_116(rr_data[115]),
                   .rr_data_117(rr_data[116]),
                   .rr_data_118(rr_data[117]),
                   .rr_data_119(rr_data[118]),
                   .rr_data_120(rr_data[119]),
                   .rr_data_121(rr_data[120]),
                   .rr_data_122(rr_data[121]),
                   .rr_data_123(rr_data[122]),
                   .rr_data_124(rr_data[123]),
                   .rr_data_125(rr_data[124]),
                   .rr_data_126(rr_data[125]),
                   .rr_data_127(rr_data[126]),
                   .rr_data_128(rr_data[127]),
                   .rr_data_129(rr_data[128]),
                   .rr_data_130(rr_data[129]),
                   .rr_data_131(rr_data[130]),
                   .rr_data_132(rr_data[131]),
                   .rr_data_133(rr_data[132]),
                   .rr_data_134(rr_data[133]),
                   .rr_data_135(rr_data[134]),
                   .rr_data_136(rr_data[135]),
                   .rr_data_137(rr_data[136]),
                   .rr_data_138(rr_data[137]),
                   .rr_data_139(rr_data[138]),
                   .rr_data_140(rr_data[139]),
                   .rr_data_141(rr_data[140]),
                   .rr_data_142(rr_data[141]),
                   .rr_data_143(rr_data[142]),
                   .rr_data_144(rr_data[143]),
                   .rr_data_145(rr_data[144]),
                   .rr_data_146(rr_data[145]),
                   .rr_data_147(rr_data[146]),
                   .rr_data_148(rr_data[147]),
                   .rr_data_149(rr_data[148]),
                   .rr_data_150(rr_data[149]),
                   .rr_data_151(rr_data[150]),
                   .rr_data_152(rr_data[151]),
                   .rr_data_153(rr_data[152]),
                   .rr_data_154(rr_data[153]),
                   .rr_data_155(rr_data[154]),
                   .rr_data_156(rr_data[155]),
                   .rr_data_157(rr_data[156]),
                   .rr_data_158(rr_data[157]),
                   .rr_data_159(rr_data[158]),
                   .rr_data_160(rr_data[159]),
                   .rr_data_161(rr_data[160]),
                   .rr_data_162(rr_data[161]),
                   .rr_data_163(rr_data[162]),
                   .rr_data_164(rr_data[163]),
                   .rr_data_165(rr_data[164]),
                   .rr_data_166(rr_data[165]),
                   .rr_data_167(rr_data[166]),
                   .rr_data_168(rr_data[167]),
                   .rr_data_169(rr_data[168]),
                   .rr_data_170(rr_data[169]),
                   .rr_data_171(rr_data[170]),
                   .rr_data_172(rr_data[171]),
                   .rr_data_173(rr_data[172]),
                   .rr_data_174(rr_data[173]),
                   .rr_data_175(rr_data[174]),
                   .rr_data_176(rr_data[175]),
                   .rr_data_177(rr_data[176]),
                   .rr_data_178(rr_data[177]),
                   .rr_data_179(rr_data[178]),
                   .rr_data_180(rr_data[179]),
                   .rr_data_181(rr_data[180]),
                   .rr_data_182(rr_data[181]),
                   .rr_data_183(rr_data[182]),
                   .rr_data_184(rr_data[183]),
                   .rr_data_185(rr_data[184]),
                   .rr_data_186(rr_data[185]),
                   .rr_data_187(rr_data[186]),
                   .rr_data_188(rr_data[187]),
                   .rr_data_189(rr_data[188]),
                   .rr_data_190(rr_data[189]),
                   .rr_data_191(rr_data[190]),
                   .rr_data_192(rr_data[191]),
                   .rr_data_193(rr_data[192]),
                   .rr_data_194(rr_data[193]),
                   .rr_data_195(rr_data[194]),
                   .rr_data_196(rr_data[195]),
                   .rr_data_197(rr_data[196]),
                   .rr_data_198(rr_data[197]),
                   .rr_data_199(rr_data[198]),
                   .rr_data_200(rr_data[199]),
                   .rr_data_201(rr_data[200]),
                   .rr_data_202(rr_data[201]),
                   .rr_data_203(rr_data[202]),
                   .rr_data_204(rr_data[203]),
                   .rr_data_205(rr_data[204]),
                   .rr_data_206(rr_data[205]),
                   .rr_data_207(rr_data[206]),
                   .rr_data_208(rr_data[207]),
                   .rr_data_209(rr_data[208]),
                   .rr_data_210(rr_data[209]),
                   .rr_data_211(rr_data[210]),
                   .rr_data_212(rr_data[211]),
                   .rr_data_213(rr_data[212]),
                   .rr_data_214(rr_data[213]),
                   .rr_data_215(rr_data[214]),
                   .rr_data_216(rr_data[215]),
                   .rr_data_217(rr_data[216]),
                   .rr_data_218(rr_data[217]),
                   .rr_data_219(rr_data[218]),
                   .rr_data_220(rr_data[219]),
                   .rr_data_221(rr_data[220]),
                   .rr_data_222(rr_data[221]),
                   .rr_data_223(rr_data[222]),
                   .rr_data_224(rr_data[223]),
                   .rr_data_225(rr_data[224]),
                   .rr_data_226(rr_data[225]),
                   .rr_data_227(rr_data[226]),
                   .rr_data_228(rr_data[227]),
                   .rr_data_229(rr_data[228]),
                   .rr_data_230(rr_data[229]),
                   .rr_data_231(rr_data[230]),
                   .rr_data_232(rr_data[231]),
                   .rr_data_233(rr_data[232]),
                   .rr_data_234(rr_data[233]),
                   .rr_data_235(rr_data[234]),
                   .rr_data_236(rr_data[235]),
                   .rr_data_237(rr_data[236]),
                   .rr_data_238(rr_data[237]),
                   .rr_data_239(rr_data[238]),
                   .rr_data_240(rr_data[239]),
                   .rr_data_241(rr_data[240]),
                   .rr_data_242(rr_data[241]),
                   .rr_data_243(rr_data[242]),
                   .rr_data_244(rr_data[243]),
                   .rr_data_245(rr_data[244]),
                   .rr_data_246(rr_data[245]),
                   .rr_data_247(rr_data[246]),
                   .rr_data_248(rr_data[247]),
                   .rr_data_249(rr_data[248]),
                   .rr_data_250(rr_data[249]),
                   .rr_data_251(rr_data[250]),
                   .rr_data_252(rr_data[251]),
                   .rr_data_253(rr_data[252]),
                   .rr_data_254(rr_data[253]),
                   .rr_data_255(rr_data[254]),
                   .rr_data_256(rr_data[255]),
                   .rr_data_257(rr_data[256]),
                   .rr_data_258(rr_data[257]),
                   .rr_data_259(rr_data[258]),
                   .rr_data_260(rr_data[259]),
                   .rr_data_261(rr_data[260]),
                   .rr_data_262(rr_data[261]),
                   .rr_data_263(rr_data[262]),
                   .rr_data_264(rr_data[263]),
                   .rr_data_265(rr_data[264]),
                   .rr_data_266(rr_data[265]),
                   .rr_data_267(rr_data[266]),
                   .rr_data_268(rr_data[267]),
                   .rr_data_269(rr_data[268]),
                   .rr_data_270(rr_data[269]),
                   .rr_data_271(rr_data[270]),
                   .rr_data_272(rr_data[271]),
                   .rr_data_273(rr_data[272]),
                   .rr_data_274(rr_data[273]),
                   .rr_data_275(rr_data[274]),
                   .rr_data_276(rr_data[275]),
                   .rr_data_277(rr_data[276]),
                   .rr_data_278(rr_data[277]),
                   .rr_data_279(rr_data[278]),
                   .rr_data_280(rr_data[279]),
                   .rr_data_281(rr_data[280]),
                   .rr_data_282(rr_data[281]),
                   .rr_data_283(rr_data[282]),
                   .rr_data_284(rr_data[283]),
                   .rr_data_285(rr_data[284]),
                   .rr_data_286(rr_data[285]),
                   .rr_data_287(rr_data[286]),
                   .rr_data_288(rr_data[287]),
                   .rr_data_289(rr_data[288]),
                   .rr_data_290(rr_data[289]),
                   .rr_data_291(rr_data[290]),
                   .rr_data_292(rr_data[291]),
                   .rr_data_293(rr_data[292]),
                   .rr_data_294(rr_data[293]),
                   .rr_data_295(rr_data[294]),
                   .rr_data_296(rr_data[295]),
                   .rr_data_297(rr_data[296]),
                   .rr_data_298(rr_data[297]),
                   .rr_data_299(rr_data[298]),
                   .rr_data_300(rr_data[299]),
                   .rr_data_301(rr_data[300]),
                   .rr_data_302(rr_data[301]),
                   .rr_data_303(rr_data[302]),
                   .rr_data_304(rr_data[303]),
                   .rr_data_305(rr_data[304]),
                   .rr_data_306(rr_data[305]),
                   .rr_data_307(rr_data[306]),
                   .rr_data_308(rr_data[307]),
                   .rr_data_309(rr_data[308]),
                   .rr_data_310(rr_data[309]),
                   .rr_data_311(rr_data[310]),
                   .rr_data_312(rr_data[311]),
                   .rr_data_313(rr_data[312]),
                   .rr_data_314(rr_data[313]),
                   .rr_data_315(rr_data[314]),
                   .rr_data_316(rr_data[315]),
                   .rr_data_317(rr_data[316]),
                   .rr_data_318(rr_data[317]),
                   .rr_data_319(rr_data[318]),
                   .rr_data_320(rr_data[319]),
                   .rr_data_321(rr_data[320]),
                   .rr_data_322(rr_data[321]),
                   .rr_data_323(rr_data[322]),
                   .rr_data_324(rr_data[323]),
                   .rr_data_325(rr_data[324]),
                   .rr_data_326(rr_data[325]),
                   .rr_data_327(rr_data[326]),
                   .rr_data_328(rr_data[327]),
                   .rr_data_329(rr_data[328]),
                   .rr_data_330(rr_data[329]),
                   .rr_data_331(rr_data[330]),
                   .rr_data_332(rr_data[331]),
                   .rr_data_333(rr_data[332]),
                   .rr_data_334(rr_data[333]),
                   .rr_data_335(rr_data[334]),
                   .rr_data_336(rr_data[335]),
                   .rr_data_337(rr_data[336]),
                   .rr_data_338(rr_data[337]),
                   .rr_data_339(rr_data[338]),
                   .rr_data_340(rr_data[339]),
                   .rr_data_341(rr_data[340]),
                   .rr_data_342(rr_data[341]),
                   .rr_data_343(rr_data[342]),
                   .rr_data_344(rr_data[343]),
                   .rr_data_345(rr_data[344]),
                   .rr_data_346(rr_data[345]),
                   .rr_data_347(rr_data[346]),
                   .rr_data_348(rr_data[347]),
                   .rr_data_349(rr_data[348]),
                   .rr_data_350(rr_data[349]),
                   .rr_data_351(rr_data[350]),
                   .rr_data_352(rr_data[351]),
                   .rr_data_353(rr_data[352]),
                   .rr_data_354(rr_data[353]),
                   .rr_data_355(rr_data[354]),
                   .rr_data_356(rr_data[355]),
                   .rr_data_357(rr_data[356]),
                   .rr_data_358(rr_data[357]),
                   .rr_data_359(rr_data[358]),
                   .rr_data_360(rr_data[359]),
                   .rr_data_361(rr_data[360]),
                   .rr_data_362(rr_data[361]),
                   .rr_data_363(rr_data[362]),
                   .rr_data_364(rr_data[363]),
                   .rr_data_365(rr_data[364]),
                   .rr_data_366(rr_data[365]),
                   .rr_data_367(rr_data[366]),
                   .rr_data_368(rr_data[367]),
                   .rr_data_369(rr_data[368]),
                   .rr_data_370(rr_data[369]),
                   .rr_data_371(rr_data[370]),
                   .rr_data_372(rr_data[371]),
                   .rr_data_373(rr_data[372]),
                   .rr_data_374(rr_data[373]),
                   .rr_data_375(rr_data[374]),
                   .rr_data_376(rr_data[375]),
                   .rr_data_377(rr_data[376]),
                   .rr_data_378(rr_data[377]),
                   .rr_data_379(rr_data[378]),
                   .rr_data_380(rr_data[379]),
                   .rr_data_381(rr_data[380]),
                   .rr_data_382(rr_data[381]),
                   .rr_data_383(rr_data[382]),
                   .rr_data_384(rr_data[383]),
                   .rr_data_385(rr_data[384]),
                   .rr_data_386(rr_data[385]),
                   .rr_data_387(rr_data[386]),
                   .rr_data_388(rr_data[387]),
                   .rr_data_389(rr_data[388]),
                   .rr_data_390(rr_data[389]),
                   .rr_data_391(rr_data[390]),
                   .rr_data_392(rr_data[391]),
                   .rr_data_393(rr_data[392]),
                   .rr_data_394(rr_data[393]),
                   .rr_data_395(rr_data[394]),
                   .rr_data_396(rr_data[395]),
                   .rr_data_397(rr_data[396]),
                   .rr_data_398(rr_data[397]),
                   .rr_data_399(rr_data[398]),
                   .rr_data_400(rr_data[399]),
                   .rr_data_401(rr_data[400]),
                   .rr_data_402(rr_data[401]),
                   .rr_data_403(rr_data[402]),
                   .rr_data_404(rr_data[403]),
                   .rr_data_405(rr_data[404]),
                   .rr_data_406(rr_data[405]),
                   .rr_data_407(rr_data[406]),
                   .rr_data_408(rr_data[407]),
                   .rr_data_409(rr_data[408]),
                   .rr_data_410(rr_data[409]),
                   .rr_data_411(rr_data[410]),
                   .rr_data_412(rr_data[411]),
                   .rr_data_413(rr_data[412]),
                   .rr_data_414(rr_data[413]),
                   .rr_data_415(rr_data[414]),
                   .rr_data_416(rr_data[415]),
                   .rr_data_417(rr_data[416]),
                   .rr_data_418(rr_data[417]),
                   .rr_data_419(rr_data[418]),
                   .rr_data_420(rr_data[419]),
                   .rr_data_421(rr_data[420]),
                   .rr_data_422(rr_data[421]),
                   .rr_data_423(rr_data[422]),
                   .rr_data_424(rr_data[423]),
                   .rr_data_425(rr_data[424]),
                   .rr_data_426(rr_data[425]),
                   .rr_data_427(rr_data[426]),
                   .rr_data_428(rr_data[427]),
                   .rr_data_429(rr_data[428]),
                   .rr_data_430(rr_data[429]),
                   .rr_data_431(rr_data[430]),
                   .rr_data_432(rr_data[431]),
                   .rr_data_433(rr_data[432]),
                   .rr_data_434(rr_data[433]),
                   .rr_data_435(rr_data[434]),
                   .rr_data_436(rr_data[435]),
                   .rr_data_437(rr_data[436]),
                   .rr_data_438(rr_data[437]),
                   .rr_data_439(rr_data[438]),
                   .rr_data_440(rr_data[439]),
                   .rr_data_441(rr_data[440]),
                   .rr_data_442(rr_data[441]),
                   .rr_data_443(rr_data[442]),
                   .rr_data_444(rr_data[443]),
                   .rr_data_445(rr_data[444]),
                   .rr_data_446(rr_data[445]),
                   .rr_data_447(rr_data[446]),
                   .rr_data_448(rr_data[447]),
                   .rr_data_449(rr_data[448]),
                   .rr_data_450(rr_data[449]),
                   .rr_data_451(rr_data[450]),
                   .rr_data_452(rr_data[451]),
                   .rr_data_453(rr_data[452]),
                   .rr_data_454(rr_data[453]),
                   .rr_data_455(rr_data[454]),
                   .rr_data_456(rr_data[455]),
                   .rr_data_457(rr_data[456]),
                   .rr_data_458(rr_data[457]),
                   .rr_data_459(rr_data[458]),
                   .rr_data_460(rr_data[459]),
                   .rr_data_461(rr_data[460]),
                   .rr_data_462(rr_data[461]),
                   .rr_data_463(rr_data[462]),
                   .rr_data_464(rr_data[463]),
                   .rr_data_465(rr_data[464]),
                   .rr_data_466(rr_data[465]),
                   .rr_data_467(rr_data[466]),
                   .rr_data_468(rr_data[467]),
                   .rr_data_469(rr_data[468]),
                   .rr_data_470(rr_data[469]),
                   .rr_data_471(rr_data[470]),
                   .rr_data_472(rr_data[471]),
                   .rr_data_473(rr_data[472]),
                   .rr_data_474(rr_data[473]),
                   .rr_data_475(rr_data[474]),
                   .rr_data_476(rr_data[475]),
                   .rr_data_477(rr_data[476]),
                   .rr_data_478(rr_data[477]),
                   .rr_data_479(rr_data[478]),
                   .rr_data_480(rr_data[479]),
                   .rr_data_481(rr_data[480]),
                   .rr_data_482(rr_data[481]),
                   .rr_data_483(rr_data[482]),
                   .rr_data_484(rr_data[483]),
                   .rr_data_485(rr_data[484]),
                   .rr_data_486(rr_data[485]),
                   .rr_data_487(rr_data[486]),
                   .rr_data_488(rr_data[487]),
                   .rr_data_489(rr_data[488]),
                   .rr_data_490(rr_data[489]),
                   .rr_data_491(rr_data[490]),
                   .rr_data_492(rr_data[491]),
                   .rr_data_493(rr_data[492]),
                   .rr_data_494(rr_data[493]),
                   .rr_data_495(rr_data[494]),
                   .rr_data_496(rr_data[495]),
                   .rr_data_497(rr_data[496]),
                   .rr_data_498(rr_data[497]),
                   .rr_data_499(rr_data[498]),
                   .rr_data_500(rr_data[499]),
                   .rr_data_501(rr_data[500]),
                   .rr_data_502(rr_data[501]),
                   .rr_data_503(rr_data[502]),
                   .rr_data_504(rr_data[503]),
                   .rr_data_505(rr_data[504]),
                   .rr_data_506(rr_data[505]),
                   .rr_data_507(rr_data[506]),
                   .rr_data_508(rr_data[507]),
                   .rr_data_509(rr_data[508]),
                   .rr_data_510(rr_data[509]),
                   .rr_data_511(rr_data[510]),
                   .rr_data_512(rr_data[511]),
                   .rr_data_513(rr_data[512]),
                   .rr_data_514(rr_data[513]),
                   .rr_data_515(rr_data[514]),
                   .rr_data_516(rr_data[515]),
                   .rr_data_517(rr_data[516]),
                   .rr_data_518(rr_data[517]),
                   .rr_data_519(rr_data[518]),
                   .rr_data_520(rr_data[519]),
                   .rr_data_521(rr_data[520]),
                   .rr_data_522(rr_data[521]),
                   .rr_data_523(rr_data[522]),
                   .rr_data_524(rr_data[523]),
                   .rr_data_525(rr_data[524]),
                   .rr_data_526(rr_data[525]),
                   .rr_data_527(rr_data[526]),
                   .rr_data_528(rr_data[527]),
                   .rr_data_529(rr_data[528]),
                   .rr_data_530(rr_data[529]),
                   .rr_data_531(rr_data[530]),
                   .rr_data_532(rr_data[531]),
                   .rr_data_533(rr_data[532]),

                  .addr          (buffer_addr),
                  .flag_buffer_in(flag_buffer_in),
                  .flag_org_write_end(flag_org_write_end),
                  .buffer_full   (buffer_full)
              );


    conctrl conctrl_inst (
                .sys_clk          (sys_clk),
                .sys_rst_n        (sys_rst_n),
                .flag_buffer_in   (flag_buffer_in),
                .flag_org_write_end(flag_org_write_end),
                .flag_org_read_end(flag_org_read_end),
                .flag_VFU_end     (flag_VFU_end),
                .flag_CFU_end     (flag_CFU_end),
                .flag_judge_end   (flag_judge_end),
                .H_sum            (H_sum),

                .flag_first_store   (flag_first_store),
                .flag_org_read_start(flag_org_read_start),
                .flag_VFU_start     (flag_VFU_start),
                .flag_CFU_start     (flag_CFU_start),
                .flag_judge_start   (flag_judge_start),
                .flag_serial        (flag_serial),
                .flag_org_update    (flag_org_update),
                .iter               (iter)
            );


    // 533 个 ram 存储输入的原始 llr 数据
`include "combine_ram_llr_1_533.txt"
    /* combine_ram_llr	combine_ram_llr_inst_1
    (
	.sys_clk		(sys_clk),
	.sys_rst_n		(sys_rst_n),
	.flag_org_read_start(flag_org_read_start),
	.buffer_addr	(buffer_addr),
	.rr_data		(rr_data[0]),
	.buffer_wr_en	(buffer_wr_en),
	.org_data		(org_data[1][15:0]),
	.org_addr		(org_addr[1][4:0]),
	.org_wr_en		(org_wr_en[1]),
	.flag_org_read_end(flag_org_read_end[0])
    ); */


    // 定义 H 扩展矩阵
`include "Hb_H_QC_N68224_K65536_R0.96_z128.txt"
    /* parameter  cyclic_shif_data_1_2   =   6'd23; */


    // 76个存储单元
`include "combine_ram_ctrl_inst21_533.txt"
    /* combine_ram_ctrl		ram_ctrl_inst_1_2 //有76个单元
    (
    .sys_clk			(sys_clk		),
    .sys_rst_n			(sys_rst_n		),
    .flag_first_store	(flag_first_store),

    .org_addr	(org_addr[2]	),
    .org_data	(org_data[2]),
    .org_wr_en	(org_wr_en[2]	),
    .VFU_addr	(VFU_addr_2	),
    .VFU_data	(VFU_data_1_2	),
    .VFU_wr_en	(VFU_wr_en_2),
    .VFU_re_en	(VFU_re_en_2),
    .cyclic_shif(cyclic_shif_data_1_2),	

    .ram_port_2_data	(CFU_data_1_2),
    .ram_port_2_wr_en	(CFU_wr_en_1),
    .ram_port_2_addr	(CFU_addr_1),
    .ram_port_2_rd_en	(CFU_re_en_1),

    .q_a_data(ram_VFU_data_1_2),
    .q_b_data(ram_CFU_data_1_2)
    ); */


    // 12个校验节点计算模块，6意味着权重行权重为6，7意味着行权重为7
`include "CFU_inst_1_21.txt"
    /* CFU_6_ctrl	CFU_6_ctrl_1
    (
    .sys_clk			(sys_clk		),
    .sys_rst_n			(sys_rst_n		),
    .flag_CFU_start	(flag_CFU_start),
    .ram_CFU_data_1	(ram_CFU_data_1_2	),//ram_port1的数据输出
    .ram_CFU_data_2	(ram_CFU_data_1_3	),//ram_port1的数据输出
    .ram_CFU_data_3	(ram_CFU_data_1_9	),//ram_port1的数据输出
    .ram_CFU_data_4	(ram_CFU_data_1_10	),//ram_port1的数据输出
    .ram_CFU_data_5	(ram_CFU_data_1_13	),//ram_port1的数据输出
    .ram_CFU_data_6	(ram_CFU_data_1_14	),//ram_port1的数据输出
    .CFU_data_7	(CFU_data_1_2	),
    .CFU_data_8	(CFU_data_1_3	),
    .CFU_data_9	(CFU_data_1_9	),
    .CFU_data_10	(CFU_data_1_10	),
    .CFU_data_11	(CFU_data_1_13	),
    .CFU_data_12	(CFU_data_1_14	),
    .CFU_addr	(CFU_addr_1	),
    .CFU_wr_en	(CFU_wr_en_1),//CFU的写使能	
    .CFU_re_en	(CFU_re_en_1),//CFU的读使能
    .flag_CFU_end	(flag_CFU_end)
    ); */


    // 24个变量节点计算模块，更新变量节点数据并计算硬判决数据
`include "VFU_inst_1_533.txt"
    /* VFU_3_ctrl	VFU_3_ctrl_1
    (
    .sys_clk		(sys_clk		),
    .sys_rst_n		(sys_rst_n		),
    .flag_VFU_start	(flag_VFU_start),
    .org_data		(org_data[1]	),
    .ram_VFU_data_1	(ram_VFU_data_4_1	),
    .ram_VFU_data_2	(ram_VFU_data_9_1	),
    .ram_VFU_data_3	(ram_VFU_data_12_1	),



    .VFU_data_1		(VFU_data_4_1	),
    .VFU_data_2		(VFU_data_9_1	),
    .VFU_data_3		(VFU_data_12_1	),
    .VFU_addr		(VFU_addr_1	),
    .VFU_wr_en		(VFU_wr_en_1),//VFU的写使能
    .VFU_re_en		(VFU_re_en_1),//VFU的读使能
    .bit_data_reg	(bit_data[0]),//硬判决数据
    .flag_VFU_end	(flag_VFU_end[0])
    ); */


    // 判决模块
    judge_ctrl judge_ctrl_inst (
                   .sys_clk         (sys_clk),
                   .sys_rst_n       (sys_rst_n),
                   .flag_judge_start(flag_judge_start),

                   .bit_data_1  (bit_data[0 ]),

                   .bit_data_2  (bit_data[1 ]),

                   .bit_data_3  (bit_data[2 ]),

                   .bit_data_4  (bit_data[3 ]),

                   .bit_data_5  (bit_data[4 ]),

                   .bit_data_6  (bit_data[5 ]),

                   .bit_data_7  (bit_data[6 ]),

                   .bit_data_8  (bit_data[7 ]),

                   .bit_data_9  (bit_data[8 ]),

                   .bit_data_10 (bit_data[9 ]),

                   .bit_data_11 (bit_data[10]),

                   .bit_data_12 (bit_data[11]),

                   .bit_data_13 (bit_data[12]),

                   .bit_data_14 (bit_data[13]),

                   .bit_data_15 (bit_data[14]),

                   .bit_data_16 (bit_data[15]),

                   .bit_data_17 (bit_data[16]),

                   .bit_data_18 (bit_data[17]),

                   .bit_data_19 (bit_data[18]),

                   .bit_data_20 (bit_data[19]),

                   .bit_data_21 (bit_data[20]),

                   .bit_data_22 (bit_data[21]),

                   .bit_data_23 (bit_data[22]),

                   .bit_data_24 (bit_data[23]),

                   .bit_data_25 (bit_data[24]),

                   .bit_data_26 (bit_data[25]),

                   .bit_data_27 (bit_data[26]),

                   .bit_data_28 (bit_data[27]),

                   .bit_data_29 (bit_data[28]),

                   .bit_data_30 (bit_data[29]),

                   .bit_data_31 (bit_data[30]),

                   .bit_data_32 (bit_data[31]),

                   .bit_data_33 (bit_data[32]),

                   .bit_data_34 (bit_data[33]),

                   .bit_data_35 (bit_data[34]),

                   .bit_data_36 (bit_data[35]),

                   .bit_data_37 (bit_data[36]),

                   .bit_data_38 (bit_data[37]),

                   .bit_data_39 (bit_data[38]),

                   .bit_data_40 (bit_data[39]),

                   .bit_data_41 (bit_data[40]),

                   .bit_data_42 (bit_data[41]),

                   .bit_data_43 (bit_data[42]),

                   .bit_data_44 (bit_data[43]),

                   .bit_data_45 (bit_data[44]),

                   .bit_data_46 (bit_data[45]),

                   .bit_data_47 (bit_data[46]),

                   .bit_data_48 (bit_data[47]),

                   .bit_data_49 (bit_data[48]),

                   .bit_data_50 (bit_data[49]),

                   .bit_data_51 (bit_data[50]),

                   .bit_data_52 (bit_data[51]),

                   .bit_data_53 (bit_data[52]),

                   .bit_data_54 (bit_data[53]),

                   .bit_data_55 (bit_data[54]),

                   .bit_data_56 (bit_data[55]),

                   .bit_data_57 (bit_data[56]),

                   .bit_data_58 (bit_data[57]),

                   .bit_data_59 (bit_data[58]),

                   .bit_data_60 (bit_data[59]),

                   .bit_data_61 (bit_data[60]),

                   .bit_data_62 (bit_data[61]),

                   .bit_data_63 (bit_data[62]),

                   .bit_data_64 (bit_data[63]),

                   .bit_data_65 (bit_data[64]),

                   .bit_data_66 (bit_data[65]),

                   .bit_data_67 (bit_data[66]),

                   .bit_data_68 (bit_data[67]),

                   .bit_data_69 (bit_data[68]),

                   .bit_data_70 (bit_data[69]),

                   .bit_data_71 (bit_data[70]),

                   .bit_data_72 (bit_data[71]),

                   .bit_data_73 (bit_data[72]),

                   .bit_data_74 (bit_data[73]),

                   .bit_data_75 (bit_data[74]),

                   .bit_data_76 (bit_data[75]),

                   .bit_data_77 (bit_data[76]),

                   .bit_data_78 (bit_data[77]),

                   .bit_data_79 (bit_data[78]),

                   .bit_data_80 (bit_data[79]),

                   .bit_data_81 (bit_data[80]),

                   .bit_data_82 (bit_data[81]),

                   .bit_data_83 (bit_data[82]),

                   .bit_data_84 (bit_data[83]),

                   .bit_data_85 (bit_data[84]),

                   .bit_data_86 (bit_data[85]),

                   .bit_data_87 (bit_data[86]),

                   .bit_data_88 (bit_data[87]),

                   .bit_data_89 (bit_data[88]),

                   .bit_data_90 (bit_data[89]),

                   .bit_data_91 (bit_data[90]),

                   .bit_data_92 (bit_data[91]),

                   .bit_data_93 (bit_data[92]),

                   .bit_data_94 (bit_data[93]),

                   .bit_data_95 (bit_data[94]),

                   .bit_data_96 (bit_data[95]),

                   .bit_data_97 (bit_data[96]),

                   .bit_data_98 (bit_data[97]),

                   .bit_data_99 (bit_data[98]),

                   .bit_data_100(bit_data[99]),

                   .bit_data_101(bit_data[100]),
                   .bit_data_102(bit_data[101]),
                   .bit_data_103(bit_data[102]),
                   .bit_data_104(bit_data[103]),
                   .bit_data_105(bit_data[104]),
                   .bit_data_106(bit_data[105]),
                   .bit_data_107(bit_data[106]),
                   .bit_data_108(bit_data[107]),
                   .bit_data_109(bit_data[108]),
                   .bit_data_110(bit_data[109]),
                   .bit_data_111(bit_data[110]),
                   .bit_data_112(bit_data[111]),
                   .bit_data_113(bit_data[112]),
                   .bit_data_114(bit_data[113]),
                   .bit_data_115(bit_data[114]),
                   .bit_data_116(bit_data[115]),
                   .bit_data_117(bit_data[116]),
                   .bit_data_118(bit_data[117]),
                   .bit_data_119(bit_data[118]),
                   .bit_data_120(bit_data[119]),
                   .bit_data_121(bit_data[120]),
                   .bit_data_122(bit_data[121]),
                   .bit_data_123(bit_data[122]),
                   .bit_data_124(bit_data[123]),
                   .bit_data_125(bit_data[124]),
                   .bit_data_126(bit_data[125]),
                   .bit_data_127(bit_data[126]),
                   .bit_data_128(bit_data[127]),
                   .bit_data_129(bit_data[128]),
                   .bit_data_130(bit_data[129]),
                   .bit_data_131(bit_data[130]),
                   .bit_data_132(bit_data[131]),
                   .bit_data_133(bit_data[132]),
                   .bit_data_134(bit_data[133]),
                   .bit_data_135(bit_data[134]),
                   .bit_data_136(bit_data[135]),
                   .bit_data_137(bit_data[136]),
                   .bit_data_138(bit_data[137]),
                   .bit_data_139(bit_data[138]),
                   .bit_data_140(bit_data[139]),
                   .bit_data_141(bit_data[140]),
                   .bit_data_142(bit_data[141]),
                   .bit_data_143(bit_data[142]),
                   .bit_data_144(bit_data[143]),
                   .bit_data_145(bit_data[144]),
                   .bit_data_146(bit_data[145]),
                   .bit_data_147(bit_data[146]),
                   .bit_data_148(bit_data[147]),
                   .bit_data_149(bit_data[148]),
                   .bit_data_150(bit_data[149]),
                   .bit_data_151(bit_data[150]),
                   .bit_data_152(bit_data[151]),
                   .bit_data_153(bit_data[152]),
                   .bit_data_154(bit_data[153]),
                   .bit_data_155(bit_data[154]),
                   .bit_data_156(bit_data[155]),
                   .bit_data_157(bit_data[156]),
                   .bit_data_158(bit_data[157]),
                   .bit_data_159(bit_data[158]),
                   .bit_data_160(bit_data[159]),
                   .bit_data_161(bit_data[160]),
                   .bit_data_162(bit_data[161]),
                   .bit_data_163(bit_data[162]),
                   .bit_data_164(bit_data[163]),
                   .bit_data_165(bit_data[164]),
                   .bit_data_166(bit_data[165]),
                   .bit_data_167(bit_data[166]),
                   .bit_data_168(bit_data[167]),
                   .bit_data_169(bit_data[168]),
                   .bit_data_170(bit_data[169]),
                   .bit_data_171(bit_data[170]),
                   .bit_data_172(bit_data[171]),
                   .bit_data_173(bit_data[172]),
                   .bit_data_174(bit_data[173]),
                   .bit_data_175(bit_data[174]),
                   .bit_data_176(bit_data[175]),
                   .bit_data_177(bit_data[176]),
                   .bit_data_178(bit_data[177]),
                   .bit_data_179(bit_data[178]),
                   .bit_data_180(bit_data[179]),
                   .bit_data_181(bit_data[180]),
                   .bit_data_182(bit_data[181]),
                   .bit_data_183(bit_data[182]),
                   .bit_data_184(bit_data[183]),
                   .bit_data_185(bit_data[184]),
                   .bit_data_186(bit_data[185]),
                   .bit_data_187(bit_data[186]),
                   .bit_data_188(bit_data[187]),
                   .bit_data_189(bit_data[188]),
                   .bit_data_190(bit_data[189]),
                   .bit_data_191(bit_data[190]),
                   .bit_data_192(bit_data[191]),
                   .bit_data_193(bit_data[192]),
                   .bit_data_194(bit_data[193]),
                   .bit_data_195(bit_data[194]),
                   .bit_data_196(bit_data[195]),
                   .bit_data_197(bit_data[196]),
                   .bit_data_198(bit_data[197]),
                   .bit_data_199(bit_data[198]),
                   .bit_data_200(bit_data[199]),
                   .bit_data_201(bit_data[200]),
                   .bit_data_202(bit_data[201]),
                   .bit_data_203(bit_data[202]),
                   .bit_data_204(bit_data[203]),
                   .bit_data_205(bit_data[204]),
                   .bit_data_206(bit_data[205]),
                   .bit_data_207(bit_data[206]),
                   .bit_data_208(bit_data[207]),
                   .bit_data_209(bit_data[208]),
                   .bit_data_210(bit_data[209]),
                   .bit_data_211(bit_data[210]),
                   .bit_data_212(bit_data[211]),
                   .bit_data_213(bit_data[212]),
                   .bit_data_214(bit_data[213]),
                   .bit_data_215(bit_data[214]),
                   .bit_data_216(bit_data[215]),
                   .bit_data_217(bit_data[216]),
                   .bit_data_218(bit_data[217]),
                   .bit_data_219(bit_data[218]),
                   .bit_data_220(bit_data[219]),
                   .bit_data_221(bit_data[220]),
                   .bit_data_222(bit_data[221]),
                   .bit_data_223(bit_data[222]),
                   .bit_data_224(bit_data[223]),
                   .bit_data_225(bit_data[224]),
                   .bit_data_226(bit_data[225]),
                   .bit_data_227(bit_data[226]),
                   .bit_data_228(bit_data[227]),
                   .bit_data_229(bit_data[228]),
                   .bit_data_230(bit_data[229]),
                   .bit_data_231(bit_data[230]),
                   .bit_data_232(bit_data[231]),
                   .bit_data_233(bit_data[232]),
                   .bit_data_234(bit_data[233]),
                   .bit_data_235(bit_data[234]),
                   .bit_data_236(bit_data[235]),
                   .bit_data_237(bit_data[236]),
                   .bit_data_238(bit_data[237]),
                   .bit_data_239(bit_data[238]),
                   .bit_data_240(bit_data[239]),
                   .bit_data_241(bit_data[240]),
                   .bit_data_242(bit_data[241]),
                   .bit_data_243(bit_data[242]),
                   .bit_data_244(bit_data[243]),
                   .bit_data_245(bit_data[244]),
                   .bit_data_246(bit_data[245]),
                   .bit_data_247(bit_data[246]),
                   .bit_data_248(bit_data[247]),
                   .bit_data_249(bit_data[248]),
                   .bit_data_250(bit_data[249]),
                   .bit_data_251(bit_data[250]),
                   .bit_data_252(bit_data[251]),
                   .bit_data_253(bit_data[252]),
                   .bit_data_254(bit_data[253]),
                   .bit_data_255(bit_data[254]),
                   .bit_data_256(bit_data[255]),
                   .bit_data_257(bit_data[256]),
                   .bit_data_258(bit_data[257]),
                   .bit_data_259(bit_data[258]),
                   .bit_data_260(bit_data[259]),
                   .bit_data_261(bit_data[260]),
                   .bit_data_262(bit_data[261]),
                   .bit_data_263(bit_data[262]),
                   .bit_data_264(bit_data[263]),
                   .bit_data_265(bit_data[264]),
                   .bit_data_266(bit_data[265]),
                   .bit_data_267(bit_data[266]),
                   .bit_data_268(bit_data[267]),
                   .bit_data_269(bit_data[268]),
                   .bit_data_270(bit_data[269]),
                   .bit_data_271(bit_data[270]),
                   .bit_data_272(bit_data[271]),
                   .bit_data_273(bit_data[272]),
                   .bit_data_274(bit_data[273]),
                   .bit_data_275(bit_data[274]),
                   .bit_data_276(bit_data[275]),
                   .bit_data_277(bit_data[276]),
                   .bit_data_278(bit_data[277]),
                   .bit_data_279(bit_data[278]),
                   .bit_data_280(bit_data[279]),
                   .bit_data_281(bit_data[280]),
                   .bit_data_282(bit_data[281]),
                   .bit_data_283(bit_data[282]),
                   .bit_data_284(bit_data[283]),
                   .bit_data_285(bit_data[284]),
                   .bit_data_286(bit_data[285]),
                   .bit_data_287(bit_data[286]),
                   .bit_data_288(bit_data[287]),
                   .bit_data_289(bit_data[288]),
                   .bit_data_290(bit_data[289]),
                   .bit_data_291(bit_data[290]),
                   .bit_data_292(bit_data[291]),
                   .bit_data_293(bit_data[292]),
                   .bit_data_294(bit_data[293]),
                   .bit_data_295(bit_data[294]),
                   .bit_data_296(bit_data[295]),
                   .bit_data_297(bit_data[296]),
                   .bit_data_298(bit_data[297]),
                   .bit_data_299(bit_data[298]),
                   .bit_data_300(bit_data[299]),
                   .bit_data_301(bit_data[300]),
                   .bit_data_302(bit_data[301]),
                   .bit_data_303(bit_data[302]),
                   .bit_data_304(bit_data[303]),
                   .bit_data_305(bit_data[304]),
                   .bit_data_306(bit_data[305]),
                   .bit_data_307(bit_data[306]),
                   .bit_data_308(bit_data[307]),
                   .bit_data_309(bit_data[308]),
                   .bit_data_310(bit_data[309]),
                   .bit_data_311(bit_data[310]),
                   .bit_data_312(bit_data[311]),
                   .bit_data_313(bit_data[312]),
                   .bit_data_314(bit_data[313]),
                   .bit_data_315(bit_data[314]),
                   .bit_data_316(bit_data[315]),
                   .bit_data_317(bit_data[316]),
                   .bit_data_318(bit_data[317]),
                   .bit_data_319(bit_data[318]),
                   .bit_data_320(bit_data[319]),
                   .bit_data_321(bit_data[320]),
                   .bit_data_322(bit_data[321]),
                   .bit_data_323(bit_data[322]),
                   .bit_data_324(bit_data[323]),
                   .bit_data_325(bit_data[324]),
                   .bit_data_326(bit_data[325]),
                   .bit_data_327(bit_data[326]),
                   .bit_data_328(bit_data[327]),
                   .bit_data_329(bit_data[328]),
                   .bit_data_330(bit_data[329]),
                   .bit_data_331(bit_data[330]),
                   .bit_data_332(bit_data[331]),
                   .bit_data_333(bit_data[332]),
                   .bit_data_334(bit_data[333]),
                   .bit_data_335(bit_data[334]),
                   .bit_data_336(bit_data[335]),
                   .bit_data_337(bit_data[336]),
                   .bit_data_338(bit_data[337]),
                   .bit_data_339(bit_data[338]),
                   .bit_data_340(bit_data[339]),
                   .bit_data_341(bit_data[340]),
                   .bit_data_342(bit_data[341]),
                   .bit_data_343(bit_data[342]),
                   .bit_data_344(bit_data[343]),
                   .bit_data_345(bit_data[344]),
                   .bit_data_346(bit_data[345]),
                   .bit_data_347(bit_data[346]),
                   .bit_data_348(bit_data[347]),
                   .bit_data_349(bit_data[348]),
                   .bit_data_350(bit_data[349]),
                   .bit_data_351(bit_data[350]),
                   .bit_data_352(bit_data[351]),
                   .bit_data_353(bit_data[352]),
                   .bit_data_354(bit_data[353]),
                   .bit_data_355(bit_data[354]),
                   .bit_data_356(bit_data[355]),
                   .bit_data_357(bit_data[356]),
                   .bit_data_358(bit_data[357]),
                   .bit_data_359(bit_data[358]),
                   .bit_data_360(bit_data[359]),
                   .bit_data_361(bit_data[360]),
                   .bit_data_362(bit_data[361]),
                   .bit_data_363(bit_data[362]),
                   .bit_data_364(bit_data[363]),
                   .bit_data_365(bit_data[364]),
                   .bit_data_366(bit_data[365]),
                   .bit_data_367(bit_data[366]),
                   .bit_data_368(bit_data[367]),
                   .bit_data_369(bit_data[368]),
                   .bit_data_370(bit_data[369]),
                   .bit_data_371(bit_data[370]),
                   .bit_data_372(bit_data[371]),
                   .bit_data_373(bit_data[372]),
                   .bit_data_374(bit_data[373]),
                   .bit_data_375(bit_data[374]),
                   .bit_data_376(bit_data[375]),
                   .bit_data_377(bit_data[376]),
                   .bit_data_378(bit_data[377]),
                   .bit_data_379(bit_data[378]),
                   .bit_data_380(bit_data[379]),
                   .bit_data_381(bit_data[380]),
                   .bit_data_382(bit_data[381]),
                   .bit_data_383(bit_data[382]),
                   .bit_data_384(bit_data[383]),
                   .bit_data_385(bit_data[384]),
                   .bit_data_386(bit_data[385]),
                   .bit_data_387(bit_data[386]),
                   .bit_data_388(bit_data[387]),
                   .bit_data_389(bit_data[388]),
                   .bit_data_390(bit_data[389]),
                   .bit_data_391(bit_data[390]),
                   .bit_data_392(bit_data[391]),
                   .bit_data_393(bit_data[392]),
                   .bit_data_394(bit_data[393]),
                   .bit_data_395(bit_data[394]),
                   .bit_data_396(bit_data[395]),
                   .bit_data_397(bit_data[396]),
                   .bit_data_398(bit_data[397]),
                   .bit_data_399(bit_data[398]),
                   .bit_data_400(bit_data[399]),
                   .bit_data_401(bit_data[400]),
                   .bit_data_402(bit_data[401]),
                   .bit_data_403(bit_data[402]),
                   .bit_data_404(bit_data[403]),
                   .bit_data_405(bit_data[404]),
                   .bit_data_406(bit_data[405]),
                   .bit_data_407(bit_data[406]),
                   .bit_data_408(bit_data[407]),
                   .bit_data_409(bit_data[408]),
                   .bit_data_410(bit_data[409]),
                   .bit_data_411(bit_data[410]),
                   .bit_data_412(bit_data[411]),
                   .bit_data_413(bit_data[412]),
                   .bit_data_414(bit_data[413]),
                   .bit_data_415(bit_data[414]),
                   .bit_data_416(bit_data[415]),
                   .bit_data_417(bit_data[416]),
                   .bit_data_418(bit_data[417]),
                   .bit_data_419(bit_data[418]),
                   .bit_data_420(bit_data[419]),
                   .bit_data_421(bit_data[420]),
                   .bit_data_422(bit_data[421]),
                   .bit_data_423(bit_data[422]),
                   .bit_data_424(bit_data[423]),
                   .bit_data_425(bit_data[424]),
                   .bit_data_426(bit_data[425]),
                   .bit_data_427(bit_data[426]),
                   .bit_data_428(bit_data[427]),
                   .bit_data_429(bit_data[428]),
                   .bit_data_430(bit_data[429]),
                   .bit_data_431(bit_data[430]),
                   .bit_data_432(bit_data[431]),
                   .bit_data_433(bit_data[432]),
                   .bit_data_434(bit_data[433]),
                   .bit_data_435(bit_data[434]),
                   .bit_data_436(bit_data[435]),
                   .bit_data_437(bit_data[436]),
                   .bit_data_438(bit_data[437]),
                   .bit_data_439(bit_data[438]),
                   .bit_data_440(bit_data[439]),
                   .bit_data_441(bit_data[440]),
                   .bit_data_442(bit_data[441]),
                   .bit_data_443(bit_data[442]),
                   .bit_data_444(bit_data[443]),
                   .bit_data_445(bit_data[444]),
                   .bit_data_446(bit_data[445]),
                   .bit_data_447(bit_data[446]),
                   .bit_data_448(bit_data[447]),
                   .bit_data_449(bit_data[448]),
                   .bit_data_450(bit_data[449]),
                   .bit_data_451(bit_data[450]),
                   .bit_data_452(bit_data[451]),
                   .bit_data_453(bit_data[452]),
                   .bit_data_454(bit_data[453]),
                   .bit_data_455(bit_data[454]),
                   .bit_data_456(bit_data[455]),
                   .bit_data_457(bit_data[456]),
                   .bit_data_458(bit_data[457]),
                   .bit_data_459(bit_data[458]),
                   .bit_data_460(bit_data[459]),
                   .bit_data_461(bit_data[460]),
                   .bit_data_462(bit_data[461]),
                   .bit_data_463(bit_data[462]),
                   .bit_data_464(bit_data[463]),
                   .bit_data_465(bit_data[464]),
                   .bit_data_466(bit_data[465]),
                   .bit_data_467(bit_data[466]),
                   .bit_data_468(bit_data[467]),
                   .bit_data_469(bit_data[468]),
                   .bit_data_470(bit_data[469]),
                   .bit_data_471(bit_data[470]),
                   .bit_data_472(bit_data[471]),
                   .bit_data_473(bit_data[472]),
                   .bit_data_474(bit_data[473]),
                   .bit_data_475(bit_data[474]),
                   .bit_data_476(bit_data[475]),
                   .bit_data_477(bit_data[476]),
                   .bit_data_478(bit_data[477]),
                   .bit_data_479(bit_data[478]),
                   .bit_data_480(bit_data[479]),
                   .bit_data_481(bit_data[480]),
                   .bit_data_482(bit_data[481]),
                   .bit_data_483(bit_data[482]),
                   .bit_data_484(bit_data[483]),
                   .bit_data_485(bit_data[484]),
                   .bit_data_486(bit_data[485]),
                   .bit_data_487(bit_data[486]),
                   .bit_data_488(bit_data[487]),
                   .bit_data_489(bit_data[488]),
                   .bit_data_490(bit_data[489]),
                   .bit_data_491(bit_data[490]),
                   .bit_data_492(bit_data[491]),
                   .bit_data_493(bit_data[492]),
                   .bit_data_494(bit_data[493]),
                   .bit_data_495(bit_data[494]),
                   .bit_data_496(bit_data[495]),
                   .bit_data_497(bit_data[496]),
                   .bit_data_498(bit_data[497]),
                   .bit_data_499(bit_data[498]),
                   .bit_data_500(bit_data[499]),
                   .bit_data_501(bit_data[500]),
                   .bit_data_502(bit_data[501]),
                   .bit_data_503(bit_data[502]),
                   .bit_data_504(bit_data[503]),
                   .bit_data_505(bit_data[504]),
                   .bit_data_506(bit_data[505]),
                   .bit_data_507(bit_data[506]),
                   .bit_data_508(bit_data[507]),
                   .bit_data_509(bit_data[508]),
                   .bit_data_510(bit_data[509]),
                   .bit_data_511(bit_data[510]),
                   .bit_data_512(bit_data[511]),
                   .bit_data_513(bit_data[512]),
                   .bit_data_514(bit_data[513]),
                   .bit_data_515(bit_data[514]),
                   .bit_data_516(bit_data[515]),
                   .bit_data_517(bit_data[516]),
                   .bit_data_518(bit_data[517]),
                   .bit_data_519(bit_data[518]),
                   .bit_data_520(bit_data[519]),
                   .bit_data_521(bit_data[520]),
                   .bit_data_522(bit_data[521]),
                   .bit_data_523(bit_data[522]),
                   .bit_data_524(bit_data[523]),
                   .bit_data_525(bit_data[524]),
                   .bit_data_526(bit_data[525]),
                   .bit_data_527(bit_data[526]),
                   .bit_data_528(bit_data[527]),
                   .bit_data_529(bit_data[528]),
                   .bit_data_530(bit_data[529]),
                   .bit_data_531(bit_data[530]),
                   .bit_data_532(bit_data[531]),
                   .bit_data_533(bit_data[532]),


                   .flag_judge_end(flag_judge_end),
                   .H_sum         (H_sum)
               );


    // 输出buffer
    buffer_out #(
                  .QC_LDPC_COL_COUNT (533)
              ) u_buffer_out (
                   .sys_clk    (sys_clk),
                   .sys_rst_n  (sys_rst_n),
                   .flag_serial(flag_serial),

                   .bit_data_1  (bit_data[0 ]),

                   .bit_data_2  (bit_data[1 ]),

                   .bit_data_3  (bit_data[2 ]),

                   .bit_data_4  (bit_data[3 ]),

                   .bit_data_5  (bit_data[4 ]),

                   .bit_data_6  (bit_data[5 ]),

                   .bit_data_7  (bit_data[6 ]),

                   .bit_data_8  (bit_data[7 ]),

                   .bit_data_9  (bit_data[8 ]),

                   .bit_data_10 (bit_data[9 ]),

                   .bit_data_11 (bit_data[10]),

                   .bit_data_12 (bit_data[11]),

                   .bit_data_13 (bit_data[12]),

                   .bit_data_14 (bit_data[13]),

                   .bit_data_15 (bit_data[14]),

                   .bit_data_16 (bit_data[15]),

                   .bit_data_17 (bit_data[16]),

                   .bit_data_18 (bit_data[17]),

                   .bit_data_19 (bit_data[18]),

                   .bit_data_20 (bit_data[19]),

                   .bit_data_21 (bit_data[20]),

                   .bit_data_22 (bit_data[21]),

                   .bit_data_23 (bit_data[22]),

                   .bit_data_24 (bit_data[23]),

                   .bit_data_25 (bit_data[24]),

                   .bit_data_26 (bit_data[25]),

                   .bit_data_27 (bit_data[26]),

                   .bit_data_28 (bit_data[27]),

                   .bit_data_29 (bit_data[28]),

                   .bit_data_30 (bit_data[29]),

                   .bit_data_31 (bit_data[30]),

                   .bit_data_32 (bit_data[31]),

                   .bit_data_33 (bit_data[32]),

                   .bit_data_34 (bit_data[33]),

                   .bit_data_35 (bit_data[34]),

                   .bit_data_36 (bit_data[35]),

                   .bit_data_37 (bit_data[36]),

                   .bit_data_38 (bit_data[37]),

                   .bit_data_39 (bit_data[38]),

                   .bit_data_40 (bit_data[39]),

                   .bit_data_41 (bit_data[40]),

                   .bit_data_42 (bit_data[41]),

                   .bit_data_43 (bit_data[42]),

                   .bit_data_44 (bit_data[43]),

                   .bit_data_45 (bit_data[44]),

                   .bit_data_46 (bit_data[45]),

                   .bit_data_47 (bit_data[46]),

                   .bit_data_48 (bit_data[47]),

                   .bit_data_49 (bit_data[48]),

                   .bit_data_50 (bit_data[49]),

                   .bit_data_51 (bit_data[50]),

                   .bit_data_52 (bit_data[51]),

                   .bit_data_53 (bit_data[52]),

                   .bit_data_54 (bit_data[53]),

                   .bit_data_55 (bit_data[54]),

                   .bit_data_56 (bit_data[55]),

                   .bit_data_57 (bit_data[56]),

                   .bit_data_58 (bit_data[57]),

                   .bit_data_59 (bit_data[58]),

                   .bit_data_60 (bit_data[59]),

                   .bit_data_61 (bit_data[60]),

                   .bit_data_62 (bit_data[61]),

                   .bit_data_63 (bit_data[62]),

                   .bit_data_64 (bit_data[63]),

                   .bit_data_65 (bit_data[64]),

                   .bit_data_66 (bit_data[65]),

                   .bit_data_67 (bit_data[66]),

                   .bit_data_68 (bit_data[67]),

                   .bit_data_69 (bit_data[68]),

                   .bit_data_70 (bit_data[69]),

                   .bit_data_71 (bit_data[70]),

                   .bit_data_72 (bit_data[71]),

                   .bit_data_73 (bit_data[72]),

                   .bit_data_74 (bit_data[73]),

                   .bit_data_75 (bit_data[74]),

                   .bit_data_76 (bit_data[75]),

                   .bit_data_77 (bit_data[76]),

                   .bit_data_78 (bit_data[77]),

                   .bit_data_79 (bit_data[78]),

                   .bit_data_80 (bit_data[79]),

                   .bit_data_81 (bit_data[80]),

                   .bit_data_82 (bit_data[81]),

                   .bit_data_83 (bit_data[82]),

                   .bit_data_84 (bit_data[83]),

                   .bit_data_85 (bit_data[84]),

                   .bit_data_86 (bit_data[85]),

                   .bit_data_87 (bit_data[86]),

                   .bit_data_88 (bit_data[87]),

                   .bit_data_89 (bit_data[88]),

                   .bit_data_90 (bit_data[89]),

                   .bit_data_91 (bit_data[90]),

                   .bit_data_92 (bit_data[91]),

                   .bit_data_93 (bit_data[92]),

                   .bit_data_94 (bit_data[93]),

                   .bit_data_95 (bit_data[94]),

                   .bit_data_96 (bit_data[95]),

                   .bit_data_97 (bit_data[96]),

                   .bit_data_98 (bit_data[97]),

                   .bit_data_99 (bit_data[98]),

                   .bit_data_100(bit_data[99]),

                   .bit_data_101(bit_data[100]),
                   .bit_data_102(bit_data[101]),
                   .bit_data_103(bit_data[102]),
                   .bit_data_104(bit_data[103]),
                   .bit_data_105(bit_data[104]),
                   .bit_data_106(bit_data[105]),
                   .bit_data_107(bit_data[106]),
                   .bit_data_108(bit_data[107]),
                   .bit_data_109(bit_data[108]),
                   .bit_data_110(bit_data[109]),
                   .bit_data_111(bit_data[110]),
                   .bit_data_112(bit_data[111]),
                   .bit_data_113(bit_data[112]),
                   .bit_data_114(bit_data[113]),
                   .bit_data_115(bit_data[114]),
                   .bit_data_116(bit_data[115]),
                   .bit_data_117(bit_data[116]),
                   .bit_data_118(bit_data[117]),
                   .bit_data_119(bit_data[118]),
                   .bit_data_120(bit_data[119]),
                   .bit_data_121(bit_data[120]),
                   .bit_data_122(bit_data[121]),
                   .bit_data_123(bit_data[122]),
                   .bit_data_124(bit_data[123]),
                   .bit_data_125(bit_data[124]),
                   .bit_data_126(bit_data[125]),
                   .bit_data_127(bit_data[126]),
                   .bit_data_128(bit_data[127]),
                   .bit_data_129(bit_data[128]),
                   .bit_data_130(bit_data[129]),
                   .bit_data_131(bit_data[130]),
                   .bit_data_132(bit_data[131]),
                   .bit_data_133(bit_data[132]),
                   .bit_data_134(bit_data[133]),
                   .bit_data_135(bit_data[134]),
                   .bit_data_136(bit_data[135]),
                   .bit_data_137(bit_data[136]),
                   .bit_data_138(bit_data[137]),
                   .bit_data_139(bit_data[138]),
                   .bit_data_140(bit_data[139]),
                   .bit_data_141(bit_data[140]),
                   .bit_data_142(bit_data[141]),
                   .bit_data_143(bit_data[142]),
                   .bit_data_144(bit_data[143]),
                   .bit_data_145(bit_data[144]),
                   .bit_data_146(bit_data[145]),
                   .bit_data_147(bit_data[146]),
                   .bit_data_148(bit_data[147]),
                   .bit_data_149(bit_data[148]),
                   .bit_data_150(bit_data[149]),
                   .bit_data_151(bit_data[150]),
                   .bit_data_152(bit_data[151]),
                   .bit_data_153(bit_data[152]),
                   .bit_data_154(bit_data[153]),
                   .bit_data_155(bit_data[154]),
                   .bit_data_156(bit_data[155]),
                   .bit_data_157(bit_data[156]),
                   .bit_data_158(bit_data[157]),
                   .bit_data_159(bit_data[158]),
                   .bit_data_160(bit_data[159]),
                   .bit_data_161(bit_data[160]),
                   .bit_data_162(bit_data[161]),
                   .bit_data_163(bit_data[162]),
                   .bit_data_164(bit_data[163]),
                   .bit_data_165(bit_data[164]),
                   .bit_data_166(bit_data[165]),
                   .bit_data_167(bit_data[166]),
                   .bit_data_168(bit_data[167]),
                   .bit_data_169(bit_data[168]),
                   .bit_data_170(bit_data[169]),
                   .bit_data_171(bit_data[170]),
                   .bit_data_172(bit_data[171]),
                   .bit_data_173(bit_data[172]),
                   .bit_data_174(bit_data[173]),
                   .bit_data_175(bit_data[174]),
                   .bit_data_176(bit_data[175]),
                   .bit_data_177(bit_data[176]),
                   .bit_data_178(bit_data[177]),
                   .bit_data_179(bit_data[178]),
                   .bit_data_180(bit_data[179]),
                   .bit_data_181(bit_data[180]),
                   .bit_data_182(bit_data[181]),
                   .bit_data_183(bit_data[182]),
                   .bit_data_184(bit_data[183]),
                   .bit_data_185(bit_data[184]),
                   .bit_data_186(bit_data[185]),
                   .bit_data_187(bit_data[186]),
                   .bit_data_188(bit_data[187]),
                   .bit_data_189(bit_data[188]),
                   .bit_data_190(bit_data[189]),
                   .bit_data_191(bit_data[190]),
                   .bit_data_192(bit_data[191]),
                   .bit_data_193(bit_data[192]),
                   .bit_data_194(bit_data[193]),
                   .bit_data_195(bit_data[194]),
                   .bit_data_196(bit_data[195]),
                   .bit_data_197(bit_data[196]),
                   .bit_data_198(bit_data[197]),
                   .bit_data_199(bit_data[198]),
                   .bit_data_200(bit_data[199]),
                   .bit_data_201(bit_data[200]),
                   .bit_data_202(bit_data[201]),
                   .bit_data_203(bit_data[202]),
                   .bit_data_204(bit_data[203]),
                   .bit_data_205(bit_data[204]),
                   .bit_data_206(bit_data[205]),
                   .bit_data_207(bit_data[206]),
                   .bit_data_208(bit_data[207]),
                   .bit_data_209(bit_data[208]),
                   .bit_data_210(bit_data[209]),
                   .bit_data_211(bit_data[210]),
                   .bit_data_212(bit_data[211]),
                   .bit_data_213(bit_data[212]),
                   .bit_data_214(bit_data[213]),
                   .bit_data_215(bit_data[214]),
                   .bit_data_216(bit_data[215]),
                   .bit_data_217(bit_data[216]),
                   .bit_data_218(bit_data[217]),
                   .bit_data_219(bit_data[218]),
                   .bit_data_220(bit_data[219]),
                   .bit_data_221(bit_data[220]),
                   .bit_data_222(bit_data[221]),
                   .bit_data_223(bit_data[222]),
                   .bit_data_224(bit_data[223]),
                   .bit_data_225(bit_data[224]),
                   .bit_data_226(bit_data[225]),
                   .bit_data_227(bit_data[226]),
                   .bit_data_228(bit_data[227]),
                   .bit_data_229(bit_data[228]),
                   .bit_data_230(bit_data[229]),
                   .bit_data_231(bit_data[230]),
                   .bit_data_232(bit_data[231]),
                   .bit_data_233(bit_data[232]),
                   .bit_data_234(bit_data[233]),
                   .bit_data_235(bit_data[234]),
                   .bit_data_236(bit_data[235]),
                   .bit_data_237(bit_data[236]),
                   .bit_data_238(bit_data[237]),
                   .bit_data_239(bit_data[238]),
                   .bit_data_240(bit_data[239]),
                   .bit_data_241(bit_data[240]),
                   .bit_data_242(bit_data[241]),
                   .bit_data_243(bit_data[242]),
                   .bit_data_244(bit_data[243]),
                   .bit_data_245(bit_data[244]),
                   .bit_data_246(bit_data[245]),
                   .bit_data_247(bit_data[246]),
                   .bit_data_248(bit_data[247]),
                   .bit_data_249(bit_data[248]),
                   .bit_data_250(bit_data[249]),
                   .bit_data_251(bit_data[250]),
                   .bit_data_252(bit_data[251]),
                   .bit_data_253(bit_data[252]),
                   .bit_data_254(bit_data[253]),
                   .bit_data_255(bit_data[254]),
                   .bit_data_256(bit_data[255]),
                   .bit_data_257(bit_data[256]),
                   .bit_data_258(bit_data[257]),
                   .bit_data_259(bit_data[258]),
                   .bit_data_260(bit_data[259]),
                   .bit_data_261(bit_data[260]),
                   .bit_data_262(bit_data[261]),
                   .bit_data_263(bit_data[262]),
                   .bit_data_264(bit_data[263]),
                   .bit_data_265(bit_data[264]),
                   .bit_data_266(bit_data[265]),
                   .bit_data_267(bit_data[266]),
                   .bit_data_268(bit_data[267]),
                   .bit_data_269(bit_data[268]),
                   .bit_data_270(bit_data[269]),
                   .bit_data_271(bit_data[270]),
                   .bit_data_272(bit_data[271]),
                   .bit_data_273(bit_data[272]),
                   .bit_data_274(bit_data[273]),
                   .bit_data_275(bit_data[274]),
                   .bit_data_276(bit_data[275]),
                   .bit_data_277(bit_data[276]),
                   .bit_data_278(bit_data[277]),
                   .bit_data_279(bit_data[278]),
                   .bit_data_280(bit_data[279]),
                   .bit_data_281(bit_data[280]),
                   .bit_data_282(bit_data[281]),
                   .bit_data_283(bit_data[282]),
                   .bit_data_284(bit_data[283]),
                   .bit_data_285(bit_data[284]),
                   .bit_data_286(bit_data[285]),
                   .bit_data_287(bit_data[286]),
                   .bit_data_288(bit_data[287]),
                   .bit_data_289(bit_data[288]),
                   .bit_data_290(bit_data[289]),
                   .bit_data_291(bit_data[290]),
                   .bit_data_292(bit_data[291]),
                   .bit_data_293(bit_data[292]),
                   .bit_data_294(bit_data[293]),
                   .bit_data_295(bit_data[294]),
                   .bit_data_296(bit_data[295]),
                   .bit_data_297(bit_data[296]),
                   .bit_data_298(bit_data[297]),
                   .bit_data_299(bit_data[298]),
                   .bit_data_300(bit_data[299]),
                   .bit_data_301(bit_data[300]),
                   .bit_data_302(bit_data[301]),
                   .bit_data_303(bit_data[302]),
                   .bit_data_304(bit_data[303]),
                   .bit_data_305(bit_data[304]),
                   .bit_data_306(bit_data[305]),
                   .bit_data_307(bit_data[306]),
                   .bit_data_308(bit_data[307]),
                   .bit_data_309(bit_data[308]),
                   .bit_data_310(bit_data[309]),
                   .bit_data_311(bit_data[310]),
                   .bit_data_312(bit_data[311]),
                   .bit_data_313(bit_data[312]),
                   .bit_data_314(bit_data[313]),
                   .bit_data_315(bit_data[314]),
                   .bit_data_316(bit_data[315]),
                   .bit_data_317(bit_data[316]),
                   .bit_data_318(bit_data[317]),
                   .bit_data_319(bit_data[318]),
                   .bit_data_320(bit_data[319]),
                   .bit_data_321(bit_data[320]),
                   .bit_data_322(bit_data[321]),
                   .bit_data_323(bit_data[322]),
                   .bit_data_324(bit_data[323]),
                   .bit_data_325(bit_data[324]),
                   .bit_data_326(bit_data[325]),
                   .bit_data_327(bit_data[326]),
                   .bit_data_328(bit_data[327]),
                   .bit_data_329(bit_data[328]),
                   .bit_data_330(bit_data[329]),
                   .bit_data_331(bit_data[330]),
                   .bit_data_332(bit_data[331]),
                   .bit_data_333(bit_data[332]),
                   .bit_data_334(bit_data[333]),
                   .bit_data_335(bit_data[334]),
                   .bit_data_336(bit_data[335]),
                   .bit_data_337(bit_data[336]),
                   .bit_data_338(bit_data[337]),
                   .bit_data_339(bit_data[338]),
                   .bit_data_340(bit_data[339]),
                   .bit_data_341(bit_data[340]),
                   .bit_data_342(bit_data[341]),
                   .bit_data_343(bit_data[342]),
                   .bit_data_344(bit_data[343]),
                   .bit_data_345(bit_data[344]),
                   .bit_data_346(bit_data[345]),
                   .bit_data_347(bit_data[346]),
                   .bit_data_348(bit_data[347]),
                   .bit_data_349(bit_data[348]),
                   .bit_data_350(bit_data[349]),
                   .bit_data_351(bit_data[350]),
                   .bit_data_352(bit_data[351]),
                   .bit_data_353(bit_data[352]),
                   .bit_data_354(bit_data[353]),
                   .bit_data_355(bit_data[354]),
                   .bit_data_356(bit_data[355]),
                   .bit_data_357(bit_data[356]),
                   .bit_data_358(bit_data[357]),
                   .bit_data_359(bit_data[358]),
                   .bit_data_360(bit_data[359]),
                   .bit_data_361(bit_data[360]),
                   .bit_data_362(bit_data[361]),
                   .bit_data_363(bit_data[362]),
                   .bit_data_364(bit_data[363]),
                   .bit_data_365(bit_data[364]),
                   .bit_data_366(bit_data[365]),
                   .bit_data_367(bit_data[366]),
                   .bit_data_368(bit_data[367]),
                   .bit_data_369(bit_data[368]),
                   .bit_data_370(bit_data[369]),
                   .bit_data_371(bit_data[370]),
                   .bit_data_372(bit_data[371]),
                   .bit_data_373(bit_data[372]),
                   .bit_data_374(bit_data[373]),
                   .bit_data_375(bit_data[374]),
                   .bit_data_376(bit_data[375]),
                   .bit_data_377(bit_data[376]),
                   .bit_data_378(bit_data[377]),
                   .bit_data_379(bit_data[378]),
                   .bit_data_380(bit_data[379]),
                   .bit_data_381(bit_data[380]),
                   .bit_data_382(bit_data[381]),
                   .bit_data_383(bit_data[382]),
                   .bit_data_384(bit_data[383]),
                   .bit_data_385(bit_data[384]),
                   .bit_data_386(bit_data[385]),
                   .bit_data_387(bit_data[386]),
                   .bit_data_388(bit_data[387]),
                   .bit_data_389(bit_data[388]),
                   .bit_data_390(bit_data[389]),
                   .bit_data_391(bit_data[390]),
                   .bit_data_392(bit_data[391]),
                   .bit_data_393(bit_data[392]),
                   .bit_data_394(bit_data[393]),
                   .bit_data_395(bit_data[394]),
                   .bit_data_396(bit_data[395]),
                   .bit_data_397(bit_data[396]),
                   .bit_data_398(bit_data[397]),
                   .bit_data_399(bit_data[398]),
                   .bit_data_400(bit_data[399]),
                   .bit_data_401(bit_data[400]),
                   .bit_data_402(bit_data[401]),
                   .bit_data_403(bit_data[402]),
                   .bit_data_404(bit_data[403]),
                   .bit_data_405(bit_data[404]),
                   .bit_data_406(bit_data[405]),
                   .bit_data_407(bit_data[406]),
                   .bit_data_408(bit_data[407]),
                   .bit_data_409(bit_data[408]),
                   .bit_data_410(bit_data[409]),
                   .bit_data_411(bit_data[410]),
                   .bit_data_412(bit_data[411]),
                   .bit_data_413(bit_data[412]),
                   .bit_data_414(bit_data[413]),
                   .bit_data_415(bit_data[414]),
                   .bit_data_416(bit_data[415]),
                   .bit_data_417(bit_data[416]),
                   .bit_data_418(bit_data[417]),
                   .bit_data_419(bit_data[418]),
                   .bit_data_420(bit_data[419]),
                   .bit_data_421(bit_data[420]),
                   .bit_data_422(bit_data[421]),
                   .bit_data_423(bit_data[422]),
                   .bit_data_424(bit_data[423]),
                   .bit_data_425(bit_data[424]),
                   .bit_data_426(bit_data[425]),
                   .bit_data_427(bit_data[426]),
                   .bit_data_428(bit_data[427]),
                   .bit_data_429(bit_data[428]),
                   .bit_data_430(bit_data[429]),
                   .bit_data_431(bit_data[430]),
                   .bit_data_432(bit_data[431]),
                   .bit_data_433(bit_data[432]),
                   .bit_data_434(bit_data[433]),
                   .bit_data_435(bit_data[434]),
                   .bit_data_436(bit_data[435]),
                   .bit_data_437(bit_data[436]),
                   .bit_data_438(bit_data[437]),
                   .bit_data_439(bit_data[438]),
                   .bit_data_440(bit_data[439]),
                   .bit_data_441(bit_data[440]),
                   .bit_data_442(bit_data[441]),
                   .bit_data_443(bit_data[442]),
                   .bit_data_444(bit_data[443]),
                   .bit_data_445(bit_data[444]),
                   .bit_data_446(bit_data[445]),
                   .bit_data_447(bit_data[446]),
                   .bit_data_448(bit_data[447]),
                   .bit_data_449(bit_data[448]),
                   .bit_data_450(bit_data[449]),
                   .bit_data_451(bit_data[450]),
                   .bit_data_452(bit_data[451]),
                   .bit_data_453(bit_data[452]),
                   .bit_data_454(bit_data[453]),
                   .bit_data_455(bit_data[454]),
                   .bit_data_456(bit_data[455]),
                   .bit_data_457(bit_data[456]),
                   .bit_data_458(bit_data[457]),
                   .bit_data_459(bit_data[458]),
                   .bit_data_460(bit_data[459]),
                   .bit_data_461(bit_data[460]),
                   .bit_data_462(bit_data[461]),
                   .bit_data_463(bit_data[462]),
                   .bit_data_464(bit_data[463]),
                   .bit_data_465(bit_data[464]),
                   .bit_data_466(bit_data[465]),
                   .bit_data_467(bit_data[466]),
                   .bit_data_468(bit_data[467]),
                   .bit_data_469(bit_data[468]),
                   .bit_data_470(bit_data[469]),
                   .bit_data_471(bit_data[470]),
                   .bit_data_472(bit_data[471]),
                   .bit_data_473(bit_data[472]),
                   .bit_data_474(bit_data[473]),
                   .bit_data_475(bit_data[474]),
                   .bit_data_476(bit_data[475]),
                   .bit_data_477(bit_data[476]),
                   .bit_data_478(bit_data[477]),
                   .bit_data_479(bit_data[478]),
                   .bit_data_480(bit_data[479]),
                   .bit_data_481(bit_data[480]),
                   .bit_data_482(bit_data[481]),
                   .bit_data_483(bit_data[482]),
                   .bit_data_484(bit_data[483]),
                   .bit_data_485(bit_data[484]),
                   .bit_data_486(bit_data[485]),
                   .bit_data_487(bit_data[486]),
                   .bit_data_488(bit_data[487]),
                   .bit_data_489(bit_data[488]),
                   .bit_data_490(bit_data[489]),
                   .bit_data_491(bit_data[490]),
                   .bit_data_492(bit_data[491]),
                   .bit_data_493(bit_data[492]),
                   .bit_data_494(bit_data[493]),
                   .bit_data_495(bit_data[494]),
                   .bit_data_496(bit_data[495]),
                   .bit_data_497(bit_data[496]),
                   .bit_data_498(bit_data[497]),
                   .bit_data_499(bit_data[498]),
                   .bit_data_500(bit_data[499]),
                   .bit_data_501(bit_data[500]),
                   .bit_data_502(bit_data[501]),
                   .bit_data_503(bit_data[502]),
                   .bit_data_504(bit_data[503]),
                   .bit_data_505(bit_data[504]),
                   .bit_data_506(bit_data[505]),
                   .bit_data_507(bit_data[506]),
                   .bit_data_508(bit_data[507]),
                   .bit_data_509(bit_data[508]),
                   .bit_data_510(bit_data[509]),
                   .bit_data_511(bit_data[510]),
                   .bit_data_512(bit_data[511]),
                   .bit_data_513(bit_data[512]),
                   .bit_data_514(bit_data[513]),
                   .bit_data_515(bit_data[514]),
                   .bit_data_516(bit_data[515]),
                   .bit_data_517(bit_data[516]),
                   .bit_data_518(bit_data[517]),
                   .bit_data_519(bit_data[518]),
                   .bit_data_520(bit_data[519]),
                   .bit_data_521(bit_data[520]),
                   .bit_data_522(bit_data[521]),
                   .bit_data_523(bit_data[522]),
                   .bit_data_524(bit_data[523]),
                   .bit_data_525(bit_data[524]),
                   .bit_data_526(bit_data[525]),
                   .bit_data_527(bit_data[526]),
                   .bit_data_528(bit_data[527]),
                   .bit_data_529(bit_data[528]),
                   .bit_data_530(bit_data[529]),
                   .bit_data_531(bit_data[530]),
                   .bit_data_532(bit_data[531]),
                   .bit_data_533(bit_data[532]),


                   .data_decode(data_decode),
                   .data_en    (data_en)
               );




endmodule
