module min_least_102 (
    input  wire [3:0] in_data_1,
    input  wire [3:0] in_data_2,
    input  wire [3:0] in_data_3,
    input  wire [3:0] in_data_4,
    input  wire [3:0] in_data_5,
    input  wire [3:0] in_data_6,
    input  wire [3:0] in_data_7,
    input  wire [3:0] in_data_8,
    input  wire [3:0] in_data_9,
    input  wire [3:0] in_data_10,
    input  wire [3:0] in_data_11,
    input  wire [3:0] in_data_12,
    input  wire [3:0] in_data_13,
    input  wire [3:0] in_data_14,
    input  wire [3:0] in_data_15,
    input  wire [3:0] in_data_16,
    input  wire [3:0] in_data_17,
    input  wire [3:0] in_data_18,
    input  wire [3:0] in_data_19,
    input  wire [3:0] in_data_20,
    input  wire [3:0] in_data_21,
    input  wire [3:0] in_data_22,
    input  wire [3:0] in_data_23,
    input  wire [3:0] in_data_24,
    input  wire [3:0] in_data_25,
    input  wire [3:0] in_data_26,
    input  wire [3:0] in_data_27,
    input  wire [3:0] in_data_28,
    input  wire [3:0] in_data_29,
    input  wire [3:0] in_data_30,
    input  wire [3:0] in_data_31,
    input  wire [3:0] in_data_32,
    input  wire [3:0] in_data_33,
    input  wire [3:0] in_data_34,
    input  wire [3:0] in_data_35,
    input  wire [3:0] in_data_36,
    input  wire [3:0] in_data_37,
    input  wire [3:0] in_data_38,
    input  wire [3:0] in_data_39,
    input  wire [3:0] in_data_40,
    input  wire [3:0] in_data_41,
    input  wire [3:0] in_data_42,
    input  wire [3:0] in_data_43,
    input  wire [3:0] in_data_44,
    input  wire [3:0] in_data_45,
    input  wire [3:0] in_data_46,
    input  wire [3:0] in_data_47,
    input  wire [3:0] in_data_48,
    input  wire [3:0] in_data_49,
    input  wire [3:0] in_data_50,
    input  wire [3:0] in_data_51,
    input  wire [3:0] in_data_52,
    input  wire [3:0] in_data_53,
    input  wire [3:0] in_data_54,
    input  wire [3:0] in_data_55,
    input  wire [3:0] in_data_56,
    input  wire [3:0] in_data_57,
    input  wire [3:0] in_data_58,
    input  wire [3:0] in_data_59,
    input  wire [3:0] in_data_60,
    input  wire [3:0] in_data_61,
    input  wire [3:0] in_data_62,
    input  wire [3:0] in_data_63,
    input  wire [3:0] in_data_64,
    input  wire [3:0] in_data_65,
    input  wire [3:0] in_data_66,
    input  wire [3:0] in_data_67,
    input  wire [3:0] in_data_68,
    input  wire [3:0] in_data_69,
    input  wire [3:0] in_data_70,
    input  wire [3:0] in_data_71,
    input  wire [3:0] in_data_72,
    input  wire [3:0] in_data_73,
    input  wire [3:0] in_data_74,
    input  wire [3:0] in_data_75,
    input  wire [3:0] in_data_76,
    input  wire [3:0] in_data_77,
    input  wire [3:0] in_data_78,
    input  wire [3:0] in_data_79,
    input  wire [3:0] in_data_80,
    input  wire [3:0] in_data_81,
    input  wire [3:0] in_data_82,
    input  wire [3:0] in_data_83,
    input  wire [3:0] in_data_84,
    input  wire [3:0] in_data_85,
    input  wire [3:0] in_data_86,
    input  wire [3:0] in_data_87,
    input  wire [3:0] in_data_88,
    input  wire [3:0] in_data_89,
    input  wire [3:0] in_data_90,
    input  wire [3:0] in_data_91,
    input  wire [3:0] in_data_92,
    input  wire [3:0] in_data_93,
    input  wire [3:0] in_data_94,
    input  wire [3:0] in_data_95,
    input  wire [3:0] in_data_96,
    input  wire [3:0] in_data_97,
    input  wire [3:0] in_data_98,
    input  wire [3:0] in_data_99,
    input  wire [3:0] in_data_100,
    input  wire [3:0] in_data_101,
    input  wire [3:0] in_data_102,

    output reg  [3:0] out_data_1,
    output reg  [3:0] out_data_2,
    output reg  [3:0] out_data_3,
    output reg  [3:0] out_data_4,
    output reg  [3:0] out_data_5,
    output reg  [3:0] out_data_6,
    output reg  [3:0] out_data_7,
    output reg  [3:0] out_data_8,
    output reg  [3:0] out_data_9,
    output reg  [3:0] out_data_10,
    output reg  [3:0] out_data_11,
    output reg  [3:0] out_data_12,
    output reg  [3:0] out_data_13,
    output reg  [3:0] out_data_14,
    output reg  [3:0] out_data_15,
    output reg  [3:0] out_data_16,
    output reg  [3:0] out_data_17,
    output reg  [3:0] out_data_18,
    output reg  [3:0] out_data_19,
    output reg  [3:0] out_data_20,
    output reg  [3:0] out_data_21,
    output reg  [3:0] out_data_22,
    output reg  [3:0] out_data_23,
    output reg  [3:0] out_data_24,
    output reg  [3:0] out_data_25,
    output reg  [3:0] out_data_26,
    output reg  [3:0] out_data_27,
    output reg  [3:0] out_data_28,
    output reg  [3:0] out_data_29,
    output reg  [3:0] out_data_30,
    output reg  [3:0] out_data_31,
    output reg  [3:0] out_data_32,
    output reg  [3:0] out_data_33,
    output reg  [3:0] out_data_34,
    output reg  [3:0] out_data_35,
    output reg  [3:0] out_data_36,
    output reg  [3:0] out_data_37,
    output reg  [3:0] out_data_38,
    output reg  [3:0] out_data_39,
    output reg  [3:0] out_data_40,
    output reg  [3:0] out_data_41,
    output reg  [3:0] out_data_42,
    output reg  [3:0] out_data_43,
    output reg  [3:0] out_data_44,
    output reg  [3:0] out_data_45,
    output reg  [3:0] out_data_46,
    output reg  [3:0] out_data_47,
    output reg  [3:0] out_data_48,
    output reg  [3:0] out_data_49,
    output reg  [3:0] out_data_50,
    output reg  [3:0] out_data_51,
    output reg  [3:0] out_data_52,
    output reg  [3:0] out_data_53,
    output reg  [3:0] out_data_54,
    output reg  [3:0] out_data_55,
    output reg  [3:0] out_data_56,
    output reg  [3:0] out_data_57,
    output reg  [3:0] out_data_58,
    output reg  [3:0] out_data_59,
    output reg  [3:0] out_data_60,
    output reg  [3:0] out_data_61,
    output reg  [3:0] out_data_62,
    output reg  [3:0] out_data_63,
    output reg  [3:0] out_data_64,
    output reg  [3:0] out_data_65,
    output reg  [3:0] out_data_66,
    output reg  [3:0] out_data_67,
    output reg  [3:0] out_data_68,
    output reg  [3:0] out_data_69,
    output reg  [3:0] out_data_70,
    output reg  [3:0] out_data_71,
    output reg  [3:0] out_data_72,
    output reg  [3:0] out_data_73,
    output reg  [3:0] out_data_74,
    output reg  [3:0] out_data_75,
    output reg  [3:0] out_data_76,
    output reg  [3:0] out_data_77,
    output reg  [3:0] out_data_78,
    output reg  [3:0] out_data_79,
    output reg  [3:0] out_data_80,
    output reg  [3:0] out_data_81,
    output reg  [3:0] out_data_82,
    output reg  [3:0] out_data_83,
    output reg  [3:0] out_data_84,
    output reg  [3:0] out_data_85,
    output reg  [3:0] out_data_86,
    output reg  [3:0] out_data_87,
    output reg  [3:0] out_data_88,
    output reg  [3:0] out_data_89,
    output reg  [3:0] out_data_90,
    output reg  [3:0] out_data_91,
    output reg  [3:0] out_data_92,
    output reg  [3:0] out_data_93,
    output reg  [3:0] out_data_94,
    output reg  [3:0] out_data_95,
    output reg  [3:0] out_data_96,
    output reg  [3:0] out_data_97,
    output reg  [3:0] out_data_98,
    output reg  [3:0] out_data_99,
    output reg  [3:0] out_data_100,
    output reg  [3:0] out_data_101,
    output reg  [3:0] out_data_102
);

    // internal array for convenience
    wire [3:0] in_data [0:101];
    assign in_data[0]  = in_data_1;
    assign in_data[1]  = in_data_2;
    assign in_data[2]  = in_data_3;
    assign in_data[3]  = in_data_4;
    assign in_data[4]  = in_data_5;
    assign in_data[5]  = in_data_6;
    assign in_data[6]  = in_data_7;
    assign in_data[7]  = in_data_8;
    assign in_data[8]  = in_data_9;
    assign in_data[9]  = in_data_10;
    assign in_data[10] = in_data_11;
    assign in_data[11] = in_data_12;
    assign in_data[12] = in_data_13;
    assign in_data[13] = in_data_14;
    assign in_data[14] = in_data_15;
    assign in_data[15] = in_data_16;
    assign in_data[16] = in_data_17;
    assign in_data[17] = in_data_18;
    assign in_data[18] = in_data_19;
    assign in_data[19] = in_data_20;
    assign in_data[20] = in_data_21;
    assign in_data[21] = in_data_22;
 assign in_data[22] = in_data_23;
    assign in_data[23] = in_data_24;
    assign in_data[24] = in_data_25;
    assign in_data[25] = in_data_26;
    assign in_data[26] = in_data_27;
    assign in_data[27] = in_data_28;
    assign in_data[28] = in_data_29;
    assign in_data[29] = in_data_30;
    assign in_data[30] = in_data_31;
    assign in_data[31] = in_data_32;
    assign in_data[32] = in_data_33;
    assign in_data[33] = in_data_34;
    assign in_data[34] = in_data_35;
    assign in_data[35] = in_data_36;
    assign in_data[36] = in_data_37;
    assign in_data[37] = in_data_38;
    assign in_data[38] = in_data_39;
    assign in_data[39] = in_data_40;
    assign in_data[40] = in_data_41;
    assign in_data[41] = in_data_42;
    assign in_data[42] = in_data_43;
    assign in_data[43] = in_data_44;
    assign in_data[44] = in_data_45;
    assign in_data[45] = in_data_46;
    assign in_data[46] = in_data_47;
    assign in_data[47] = in_data_48;
    assign in_data[48] = in_data_49;
    assign in_data[49] = in_data_50;
    assign in_data[50] = in_data_51;
    assign in_data[51] = in_data_52;
    assign in_data[52] = in_data_53;
    assign in_data[53] = in_data_54;
    assign in_data[54] = in_data_55;
    assign in_data[55] = in_data_56;
    assign in_data[56] = in_data_57;
    assign in_data[57] = in_data_58;
    assign in_data[58] = in_data_59;
    assign in_data[59] = in_data_60;
    assign in_data[60] = in_data_61;
    assign in_data[61] = in_data_62;
    assign in_data[62] = in_data_63;
    assign in_data[63] = in_data_64;
    assign in_data[64] = in_data_65;
    assign in_data[65] = in_data_66;
    assign in_data[66] = in_data_67;
    assign in_data[67] = in_data_68;
    assign in_data[68] = in_data_69;
    assign in_data[69] = in_data_70;
    assign in_data[70] = in_data_71;
    assign in_data[71] = in_data_72;
    assign in_data[72] = in_data_73;
    assign in_data[73] = in_data_74;
    assign in_data[74] = in_data_75;
    assign in_data[75] = in_data_76;
    assign in_data[76] = in_data_77;
    assign in_data[77] = in_data_78;
    assign in_data[78] = in_data_79;
    assign in_data[79] = in_data_80;
    assign in_data[80] = in_data_81;
    assign in_data[81] = in_data_82;
    assign in_data[82] = in_data_83;
    assign in_data[83] = in_data_84;
    assign in_data[84] = in_data_85;
    assign in_data[85] = in_data_86;
    assign in_data[86] = in_data_87;
    assign in_data[87] = in_data_88;
    assign in_data[88] = in_data_89;
    assign in_data[89] = in_data_90;
    assign in_data[90] = in_data_91;
    assign in_data[91] = in_data_92;
    assign in_data[92] = in_data_93;
    assign in_data[93] = in_data_94;
    assign in_data[94] = in_data_95;
    assign in_data[95] = in_data_96;
    assign in_data[96] = in_data_97;
    assign in_data[97] = in_data_98;
    assign in_data[98] = in_data_99;
    assign in_data[99] = in_data_100;
    assign in_data[100] = in_data_101;
    assign in_data[101] = in_data_102;

    // -------------------------
    // Layer1: 102 -> 51 pairs (direct compare of slices)
    // -------------------------
    wire [2:0] l1_min [0:50];
    wire [2:0] l1_least [0:50];

    genvar gi;
    generate
        for (gi = 0; gi < 51; gi = gi + 1) begin : GEN_L1_INLINE
            assign l1_min[gi]   = (in_data[2*gi][2:0] <= in_data[2*gi+1][2:0]) ? in_data[2*gi][2:0] : in_data[2*gi+1][2:0];
            assign l1_least[gi] = (in_data[2*gi][2:0] >  in_data[2*gi+1][2:0]) ? in_data[2*gi][2:0] : in_data[2*gi+1][2:0];
        end
    endgenerate

    // -------------------------
    // Layer2: 51 -> 26 (25 pairs + 1 passthrough)
    // -------------------------
    wire [2:0] l2_min [0:25];
    wire [2:0] l2_least [0:25];

    generate
        for (gi = 0; gi < 25; gi = gi + 1) begin : GEN_L2_INLINE
            assign l2_min[gi]   = (l1_min[2*gi] <= l1_min[2*gi+1]) ? l1_min[2*gi] : l1_min[2*gi+1];
            assign l2_least[gi] = (l1_min[2*gi] >  l1_min[2*gi+1]) ? l1_min[2*gi] : l1_min[2*gi+1];
        end
    endgenerate

    assign l2_min[25]   = l1_min[50];
    assign l2_least[25] = l1_least[50];

    // -------------------------
    // Layer3: 26 -> 13 (12 pairs + 1 passthrough)
    // -------------------------
    wire [2:0] l3_min [0:12];
    wire [2:0] l3_least [0:12];

    generate
        for (gi = 0; gi < 12; gi = gi + 1) begin : GEN_L3_INLINE
            assign l3_min[gi]   = (l2_min[2*gi] <= l2_min[2*gi+1]) ? l2_min[2*gi] : l2_min[2*gi+1];
            assign l3_least[gi] = (l2_min[2*gi] >  l2_min[2*gi+1]) ? l2_min[2*gi] : l2_min[2*gi+1];
        end
    endgenerate

    assign l3_min[12]   = l2_min[25];
    assign l3_least[12] = l2_least[25];

    // -------------------------
    // Layer4: 13 -> 7 (6 pairs + 1 passthrough)
    // -------------------------
    wire [2:0] l4_min [0:6];
    wire [2:0] l4_least [0:6];

    generate
        for (gi = 0; gi < 6; gi = gi + 1) begin : GEN_L4_INLINE
            assign l4_min[gi]   = (l3_min[2*gi] <= l3_min[2*gi+1]) ? l3_min[2*gi] : l3_min[2*gi+1];
            assign l4_least[gi] = (l3_min[2*gi] >  l3_min[2*gi+1]) ? l3_min[2*gi] : l3_min[2*gi+1];
        end
    endgenerate

    assign l4_min[6]   = l3_min[12];
    assign l4_least[6] = l3_least[12];

    // -------------------------
    // Layer5: 7 -> 4 (3 pairs + 1 passthrough)
    // -------------------------
    wire [2:0] l5_min [0:3];
    wire [2:0] l5_least [0:3];

    assign l5_min[0]   = (l4_min[0] <= l4_min[1]) ? l4_min[0] : l4_min[1];
    assign l5_least[0] = (l4_min[0] >  l4_min[1]) ? l4_min[0] : l4_min[1];

    assign l5_min[1]   = (l4_min[2] <= l4_min[3]) ? l4_min[2] : l4_min[3];
    assign l5_least[1] = (l4_min[2] >  l4_min[3]) ? l4_min[2] : l4_min[3];

    assign l5_min[2]   = (l4_min[4] <= l4_min[5]) ? l4_min[4] : l4_min[5];
    assign l5_least[2] = (l4_min[4] >  l4_min[5]) ? l4_min[4] : l4_min[5];

    assign l5_min[3]   = l4_min[6];
    assign l5_least[3] = l4_least[6];

    // -------------------------
    // Layer6: 4 -> 2 (1 pair + passthrough)
    // -------------------------
    wire [2:0] l6_min [0:1];
    wire [2:0] l6_least [0:1];

    assign l6_min[0]   = (l5_min[0] <= l5_min[1]) ? l5_min[0] : l5_min[1];
    assign l6_least[0] = (l5_min[0] >  l5_min[1]) ? l5_min[0] : l5_min[1];

    assign l6_min[1]   = (l5_min[2] <= l5_min[3]) ? l5_min[2] : l5_min[3];
    assign l6_least[1] = (l5_min[2] >  l5_min[3]) ? l5_min[2] : l5_min[3];

    // -------------------------
    // Final: 2 -> 1 (global_min & semifinal_min)
    // -------------------------
    wire [2:0] global_min;
    wire [2:0] semifinal_min;

    assign global_min   = (l6_min[0] <= l6_min[1]) ? l6_min[0] : l6_min[1];
    assign semifinal_min = (l6_min[0] >  l6_min[1]) ? l6_min[0] : l6_min[1];

    // -------------------------
    // Trace-back candidates (value-based)
    // -------------------------
    localparam [2:0] MAXV = 3'h7;

    wire [2:0] cand_l6 = (l6_min[0] == global_min) ? l6_least[0] : l6_least[1];

    wire [2:0] cand_l5;
    assign cand_l5 =
        (l5_min[0] == l6_min[0] && l6_min[0] == global_min) ? l5_least[0] :
        (l5_min[1] == l6_min[0] && l6_min[0] == global_min) ? l5_least[1] :
        (l5_min[2] == l6_min[1] && l6_min[1] == global_min) ? l5_least[2] :
        (l5_min[3] == l6_min[1] && l6_min[1] == global_min) ? l5_least[3] :
        MAXV;

    wire [2:0] cand_l4;
    assign cand_l4 =
        (l4_min[0]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l4_least[0] :
        (l4_min[1]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l4_least[1] :
        (l4_min[2]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l4_least[2] :
        (l4_min[3]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l4_least[3] :
        (l4_min[4]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l4_least[4] :
        (l4_min[5]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l4_least[5] :
        (l4_min[6]==l5_min[3] && l5_min[3]==l6_min[1] && l6_min[1]==global_min) ? l4_least[6] :
        MAXV;

    wire [2:0] cand_l3;
    assign cand_l3 =
        (l3_min[0]==l4_min[0] && l4_min[0]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l3_least[0] :
        (l3_min[1]==l4_min[0] && l4_min[0]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l3_least[1] :
        (l3_min[2]==l4_min[1] && l4_min[1]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l3_least[2] :
        (l3_min[3]==l4_min[1] && l4_min[1]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l3_least[3] :
        (l3_min[4]==l4_min[2] && l4_min[2]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l3_least[4] :
        (l3_min[5]==l4_min[2] && l4_min[2]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l3_least[5] :
        (l3_min[6]==l4_min[3] && l4_min[3]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l3_least[6] :
        (l3_min[7]==l4_min[3] && l4_min[3]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l3_least[7] :
        (l3_min[8]==l4_min[4] && l4_min[4]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l3_least[8] :
        (l3_min[9]==l4_min[4] && l4_min[4]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l3_least[9] :
        (l3_min[10]==l4_min[5] && l4_min[5]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l3_least[10] :
        (l3_min[11]==l4_min[5] && l4_min[5]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l3_least[11] :
        (l3_min[12]==l4_min[6] && l4_min[6]==l5_min[3] && l5_min[3]==l6_min[1] && l6_min[1]==global_min) ? l3_least[12] :
        MAXV;

    wire [2:0] cand_l2;
    assign cand_l2 =
        (l2_min[0]==l3_min[0] && l3_min[0]==l4_min[0] && l4_min[0]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l2_least[0] :
        (l2_min[1]==l3_min[0] && l3_min[0]==l4_min[0] && l4_min[0]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l2_least[1] :
        (l2_min[2]==l3_min[1] && l3_min[1]==l4_min[0] && l4_min[0]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l2_least[2] :
        (l2_min[3]==l3_min[1] && l3_min[1]==l4_min[0] && l4_min[0]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l2_least[3] :
        (l2_min[4]==l3_min[2] && l3_min[2]==l4_min[1] && l4_min[1]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l2_least[4] :
        (l2_min[5]==l3_min[2] && l3_min[2]==l4_min[1] && l4_min[1]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l2_least[5] :
        (l2_min[6]==l3_min[3] && l3_min[3]==l4_min[1] && l4_min[1]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l2_least[6] :
        (l2_min[7]==l3_min[3] && l3_min[3]==l4_min[1] && l4_min[1]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l2_least[7] :
        (l2_min[8]==l3_min[4] && l3_min[4]==l4_min[2] && l4_min[2]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l2_least[8] :
        (l2_min[9]==l3_min[4] && l3_min[4]==l4_min[2] && l4_min[2]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l2_least[9] :
        (l2_min[10]==l3_min[5] && l3_min[5]==l4_min[2] && l4_min[2]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l2_least[10] :
        (l2_min[11]==l3_min[5] && l3_min[5]==l4_min[2] && l4_min[2]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l2_least[11] :
        (l2_min[12]==l3_min[6] && l3_min[6]==l4_min[3] && l4_min[3]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l2_least[12] :
        (l2_min[13]==l3_min[6] && l3_min[6]==l4_min[3] && l4_min[3]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l2_least[13] :
        (l2_min[14]==l3_min[7] && l3_min[7]==l4_min[3] && l4_min[3]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l2_least[14] :
        (l2_min[15]==l3_min[7] && l3_min[7]==l4_min[3] && l4_min[3]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l2_least[15] :
        (l2_min[16]==l3_min[8] && l3_min[8]==l4_min[4] && l4_min[4]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l2_least[16] :
        (l2_min[17]==l3_min[8] && l3_min[8]==l4_min[4] && l4_min[4]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l2_least[17] :
        (l2_min[18]==l3_min[9] && l3_min[9]==l4_min[4] && l4_min[4]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l2_least[18] :
        (l2_min[19]==l3_min[9] && l3_min[9]==l4_min[4] && l4_min[4]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l2_least[19] :
        (l2_min[20]==l3_min[10] && l3_min[10]==l4_min[5] && l4_min[5]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l2_least[20] :
        (l2_min[21]==l3_min[10] && l3_min[10]==l4_min[5] && l4_min[5]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l2_least[21] :
        (l2_min[22]==l3_min[11] && l3_min[11]==l4_min[5] && l4_min[5]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l2_least[22] :
        (l2_min[23]==l3_min[11] && l3_min[11]==l4_min[5] && l4_min[5]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l2_least[23] :
        (l2_min[24]==l3_min[12] && l3_min[12]==l4_min[6] && l4_min[6]==l5_min[3] && l5_min[3]==l6_min[1] && l6_min[1]==global_min) ? l2_least[24] :
        (l2_min[25]==l3_min[12] && l3_min[12]==l4_min[6] && l4_min[6]==l5_min[3] && l5_min[3]==l6_min[1] && l6_min[1]==global_min) ? l2_least[25] :
        MAXV;

    wire [2:0] cand_l1;
    assign cand_l1 =
        (l1_min[0]==l2_min[0] && l2_min[0]==l3_min[0] && l3_min[0]==l4_min[0] && l4_min[0]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l1_least[0] :
        (l1_min[1]==l2_min[0] && l2_min[0]==l3_min[0] && l3_min[0]==l4_min[0] && l4_min[0]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l1_least[1] :
        (l1_min[2]==l2_min[1] && l2_min[1]==l3_min[0] && l3_min[0]==l4_min[0] && l4_min[0]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l1_least[2] :
        (l1_min[3]==l2_min[1] && l2_min[1]==l3_min[0] && l3_min[0]==l4_min[0] && l4_min[0]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l1_least[3] :
        (l1_min[4]==l2_min[2] && l2_min[2]==l3_min[1] && l3_min[1]==l4_min[0] && l4_min[0]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l1_least[4] :
        (l1_min[5]==l2_min[2] && l2_min[2]==l3_min[1] && l3_min[1]==l4_min[0] && l4_min[0]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l1_least[5] :
        (l1_min[6]==l2_min[3] && l2_min[3]==l3_min[1] && l3_min[1]==l4_min[0] && l4_min[0]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l1_least[6] :
        (l1_min[7]==l2_min[3] && l2_min[3]==l3_min[1] && l3_min[1]==l4_min[0] && l4_min[0]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l1_least[7] :
        (l1_min[8]==l2_min[4] && l2_min[4]==l3_min[2] && l3_min[2]==l4_min[1] && l4_min[1]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l1_least[8] :
        (l1_min[9]==l2_min[4] && l2_min[4]==l3_min[2] && l3_min[2]==l4_min[1] && l4_min[1]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l1_least[9] :
        (l1_min[10]==l2_min[5] && l2_min[5]==l3_min[2] && l3_min[2]==l4_min[1] && l4_min[1]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l1_least[10] :
        (l1_min[11]==l2_min[5] && l2_min[5]==l3_min[2] && l3_min[2]==l4_min[1] && l4_min[1]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l1_least[11] :
        (l1_min[12]==l2_min[6] && l2_min[6]==l3_min[3] && l3_min[3]==l4_min[1] && l4_min[1]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l1_least[12] :
        (l1_min[13]==l2_min[6] && l2_min[6]==l3_min[3] && l3_min[3]==l4_min[1] && l4_min[1]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l1_least[13] :
        (l1_min[14]==l2_min[7] && l2_min[7]==l3_min[3] && l3_min[3]==l4_min[1] && l4_min[1]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l1_least[14] :
        (l1_min[15]==l2_min[7] && l2_min[7]==l3_min[3] && l3_min[3]==l4_min[1] && l4_min[1]==l5_min[0] && l5_min[0]==l6_min[0] && l6_min[0]==global_min) ? l1_least[15] :
        (l1_min[16]==l2_min[8] && l2_min[8]==l3_min[4] && l3_min[4]==l4_min[2] && l4_min[2]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l1_least[16] :
        (l1_min[17]==l2_min[8] && l2_min[8]==l3_min[4] && l3_min[4]==l4_min[2] && l4_min[2]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l1_least[17] :
        (l1_min[18]==l2_min[9] && l2_min[9]==l3_min[4] && l3_min[4]==l4_min[2] && l4_min[2]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l1_least[18] :
        (l1_min[19]==l2_min[9] && l2_min[9]==l3_min[4] && l3_min[4]==l4_min[2] && l4_min[2]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l1_least[19] :
        (l1_min[20]==l2_min[10] && l2_min[10]==l3_min[5] && l3_min[5]==l4_min[2] && l4_min[2]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l1_least[20] :
        (l1_min[21]==l2_min[10] && l2_min[10]==l3_min[5] && l3_min[5]==l4_min[2] && l4_min[2]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l1_least[21] :
        (l1_min[22]==l2_min[11] && l2_min[11]==l3_min[5] && l3_min[5]==l4_min[2] && l4_min[2]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l1_least[22] :
        (l1_min[23]==l2_min[11] && l2_min[11]==l3_min[5] && l3_min[5]==l4_min[2] && l4_min[2]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l1_least[23] :
        (l1_min[24]==l2_min[12] && l2_min[12]==l3_min[6] && l3_min[6]==l4_min[3] && l4_min[3]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l1_least[24] :
        (l1_min[25]==l2_min[12] && l2_min[12]==l3_min[6] && l3_min[6]==l4_min[3] && l4_min[3]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l1_least[25] :
        (l1_min[26]==l2_min[13] && l2_min[13]==l3_min[6] && l3_min[6]==l4_min[3] && l4_min[3]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l1_least[26] :
        (l1_min[27]==l2_min[13] && l2_min[13]==l3_min[6] && l3_min[6]==l4_min[3] && l4_min[3]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l1_least[27] :
        (l1_min[28]==l2_min[14] && l2_min[14]==l3_min[7] && l3_min[7]==l4_min[3] && l4_min[3]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l1_least[28] :
        (l1_min[29]==l2_min[14] && l2_min[14]==l3_min[7] && l3_min[7]==l4_min[3] && l4_min[3]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l1_least[29] :
        (l1_min[30]==l2_min[15] && l2_min[15]==l3_min[7] && l3_min[7]==l4_min[3] && l4_min[3]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l1_least[30] :
        (l1_min[31]==l2_min[15] && l2_min[15]==l3_min[7] && l3_min[7]==l4_min[3] && l4_min[3]==l5_min[1] && l5_min[1]==l6_min[0] && l6_min[0]==global_min) ? l1_least[31] :
        (l1_min[32]==l2_min[16] && l2_min[16]==l3_min[8] && l3_min[8]==l4_min[4] && l4_min[4]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l1_least[32] :
        (l1_min[33]==l2_min[16] && l2_min[16]==l3_min[8] && l3_min[8]==l4_min[4] && l4_min[4]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l1_least[33] :
        (l1_min[34]==l2_min[17] && l2_min[17]==l3_min[8] && l3_min[8]==l4_min[4] && l4_min[4]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l1_least[34] :
        (l1_min[35]==l2_min[17] && l2_min[17]==l3_min[8] && l3_min[8]==l4_min[4] && l4_min[4]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l1_least[35] :
        (l1_min[36]==l2_min[18] && l2_min[18]==l3_min[9] && l3_min[9]==l4_min[4] && l4_min[4]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l1_least[36] :
        (l1_min[37]==l2_min[18] && l2_min[18]==l3_min[9] && l3_min[9]==l4_min[4] && l4_min[4]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l1_least[37] :
        (l1_min[38]==l2_min[19] && l2_min[19]==l3_min[9] && l3_min[9]==l4_min[4] && l4_min[4]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l1_least[38] :
        (l1_min[39]==l2_min[19] && l2_min[19]==l3_min[9] && l3_min[9]==l4_min[4] && l4_min[4]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l1_least[39] :
        (l1_min[40]==l2_min[20] && l2_min[20]==l3_min[10] && l3_min[10]==l4_min[5] && l4_min[5]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l1_least[40] :
        (l1_min[41]==l2_min[20] && l2_min[20]==l3_min[10] && l3_min[10]==l4_min[5] && l4_min[5]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l1_least[41] :
        (l1_min[42]==l2_min[21] && l2_min[21]==l3_min[10] && l3_min[10]==l4_min[5] && l4_min[5]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l1_least[42] :
        (l1_min[43]==l2_min[21] && l2_min[21]==l3_min[10] && l3_min[10]==l4_min[5] && l4_min[5]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l1_least[43] :
        (l1_min[44]==l2_min[22] && l2_min[22]==l3_min[11] && l3_min[11]==l4_min[5] && l4_min[5]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l1_least[44] :
        (l1_min[45]==l2_min[22] && l2_min[22]==l3_min[11] && l3_min[11]==l4_min[5] && l4_min[5]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l1_least[45] :
        (l1_min[46]==l2_min[23] && l2_min[23]==l3_min[11] && l3_min[11]==l4_min[5] && l4_min[5]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l1_least[46] :
        (l1_min[47]==l2_min[23] && l2_min[23]==l3_min[11] && l3_min[11]==l4_min[5] && l4_min[5]==l5_min[2] && l5_min[2]==l6_min[1] && l6_min[1]==global_min) ? l1_least[47] :
        (l1_min[48]==l2_min[24] && l2_min[24]==l3_min[12] && l3_min[12]==l4_min[6] && l4_min[6]==l5_min[3] && l5_min[3]==l6_min[1] && l6_min[1]==global_min) ? l1_least[48] :
        (l1_min[49]==l2_min[24] && l2_min[24]==l3_min[12] && l3_min[12]==l4_min[6] && l4_min[6]==l5_min[3] && l5_min[3]==l6_min[1] && l6_min[1]==global_min) ? l1_least[49] :
        (l1_min[50]==l2_min[25] && l2_min[25]==l3_min[12] && l3_min[12]==l4_min[6] && l4_min[6]==l5_min[3] && l5_min[3]==l6_min[1] && l6_min[1]==global_min) ? l1_least[50] :
        MAXV;

    wire [2:0] tmp0 = (semifinal_min < cand_l6) ? semifinal_min : cand_l6;
    wire [2:0] tmp1 = (tmp0 < cand_l5) ? tmp0 : cand_l5;
    wire [2:0] tmp2 = (tmp1 < cand_l4) ? tmp1 : cand_l4;
    wire [2:0] tmp3 = (tmp2 < cand_l3) ? tmp2 : cand_l3;
    wire [2:0] tmp4 = (tmp3 < cand_l2) ? tmp3 : cand_l2;
    wire [2:0] global_second = (tmp4 < cand_l1) ? tmp4 : cand_l1;

    // -------------------------
    // sign: XOR of all input sign bits (1-bit)
    // -------------------------
    wire sign;
    assign sign = in_data[0][3] ^ in_data[1][3] ^ in_data[2][3] ^ in_data[3][3] ^
                  in_data[4][3] ^ in_data[5][3] ^ in_data[6][3] ^ in_data[7][3] ^
                  in_data[8][3] ^ in_data[9][3] ^ in_data[10][3] ^ in_data[11][3] ^
                  in_data[12][3] ^ in_data[13][3] ^ in_data[14][3] ^ in_data[15][3] ^
                  in_data[16][3] ^ in_data[17][3] ^ in_data[18][3] ^ in_data[19][3] ^
                  in_data[20][3] ^ in_data[21][3] ^ in_data[22][3] ^ in_data[23][3] ^
                  in_data[24][3] ^ in_data[25][3] ^ in_data[26][3] ^ in_data[27][3] ^
                  in_data[28][3] ^ in_data[29][3] ^ in_data[30][3] ^ in_data[31][3] ^
                  in_data[32][3] ^ in_data[33][3] ^ in_data[34][3] ^ in_data[35][3] ^
                  in_data[36][3] ^ in_data[37][3] ^ in_data[38][3] ^ in_data[39][3] ^
                  in_data[40][3] ^ in_data[41][3] ^ in_data[42][3] ^ in_data[43][3] ^
                  in_data[44][3] ^ in_data[45][3] ^ in_data[46][3] ^ in_data[47][3] ^
                  in_data[48][3] ^ in_data[49][3] ^ in_data[50][3] ^ in_data[51][3] ^
                  in_data[52][3] ^ in_data[53][3] ^ in_data[54][3] ^ in_data[55][3] ^
                  in_data[56][3] ^ in_data[57][3] ^ in_data[58][3] ^ in_data[59][3] ^
                  in_data[60][3] ^ in_data[61][3] ^ in_data[62][3] ^ in_data[63][3] ^
                  in_data[64][3] ^ in_data[65][3] ^ in_data[66][3] ^ in_data[67][3] ^
                  in_data[68][3] ^ in_data[69][3] ^ in_data[70][3] ^ in_data[71][3] ^
                  in_data[72][3] ^ in_data[73][3] ^ in_data[74][3] ^ in_data[75][3] ^
                  in_data[76][3] ^ in_data[77][3] ^ in_data[78][3] ^ in_data[79][3] ^
                  in_data[80][3] ^ in_data[81][3] ^ in_data[82][3] ^ in_data[83][3] ^
                  in_data[84][3] ^ in_data[85][3] ^ in_data[86][3] ^ in_data[87][3] ^
                  in_data[88][3] ^ in_data[89][3] ^ in_data[90][3] ^ in_data[91][3] ^
                  in_data[92][3] ^ in_data[93][3] ^ in_data[94][3] ^ in_data[95][3] ^
                  in_data[96][3] ^ in_data[97][3] ^ in_data[98][3] ^ in_data[99][3] ^
                  in_data[100][3] ^ in_data[101][3];

    // -------------------------
    // final outputs (combinational)
    // -------------------------
    always @(*) begin
        out_data_1  = (in_data_1[2:0]  == global_min) ? {(in_data_1[3]  ^ sign), global_second} : {(in_data_1[3]  ^ sign), global_min};
        out_data_2  = (in_data_2[2:0]  == global_min) ? {(in_data_2[3]  ^ sign), global_second} : {(in_data_2[3]  ^ sign), global_min};
        out_data_3  = (in_data_3[2:0]  == global_min) ? {(in_data_3[3]  ^ sign), global_second} : {(in_data_3[3]  ^ sign), global_min};
        out_data_4  = (in_data_4[2:0]  == global_min) ? {(in_data_4[3]  ^ sign), global_second} : {(in_data_4[3]  ^ sign), global_min};
        out_data_5  = (in_data_5[2:0]  == global_min) ? {(in_data_5[3]  ^ sign), global_second} : {(in_data_5[3]  ^ sign), global_min};
        out_data_6  = (in_data_6[2:0]  == global_min) ? {(in_data_6[3]  ^ sign), global_second} : {(in_data_6[3]  ^ sign), global_min};
        out_data_7  = (in_data_7[2:0]  == global_min) ? {(in_data_7[3]  ^ sign), global_second} : {(in_data_7[3]  ^ sign), global_min};
        out_data_8  = (in_data_8[2:0]  == global_min) ? {(in_data_8[3]  ^ sign), global_second} : {(in_data_8[3]  ^ sign), global_min};
        out_data_9  = (in_data_9[2:0]  == global_min) ? {(in_data_9[3]  ^ sign), global_second} : {(in_data_9[3]  ^ sign), global_min};
        out_data_10 = (in_data_10[2:0] == global_min) ? {(in_data_10[3] ^ sign), global_second} : {(in_data_10[3] ^ sign), global_min};
        out_data_11 = (in_data_11[2:0] == global_min) ? {(in_data_11[3] ^ sign), global_second} : {(in_data_11[3] ^ sign), global_min};
        out_data_12 = (in_data_12[2:0] == global_min) ? {(in_data_12[3] ^ sign), global_second} : {(in_data_12[3] ^ sign), global_min};
        out_data_13 = (in_data_13[2:0] == global_min) ? {(in_data_13[3] ^ sign), global_second} : {(in_data_13[3] ^ sign), global_min};
        out_data_14 = (in_data_14[2:0] == global_min) ? {(in_data_14[3] ^ sign), global_second} : {(in_data_14[3] ^ sign), global_min};
        out_data_15 = (in_data_15[2:0] == global_min) ? {(in_data_15[3] ^ sign), global_second} : {(in_data_15[3] ^ sign), global_min};
        out_data_16 = (in_data_16[2:0] == global_min) ? {(in_data_16[3] ^ sign), global_second} : {(in_data_16[3] ^ sign), global_min};
        out_data_17 = (in_data_17[2:0] == global_min) ? {(in_data_17[3] ^ sign), global_second} : {(in_data_17[3] ^ sign), global_min};
        out_data_18 = (in_data_18[2:0] == global_min) ? {(in_data_18[3] ^ sign), global_second} : {(in_data_18[3] ^ sign), global_min};
        out_data_19 = (in_data_19[2:0] == global_min) ? {(in_data_19[3] ^ sign), global_second} : {(in_data_19[3] ^ sign), global_min};
        out_data_20 = (in_data_20[2:0] == global_min) ? {(in_data_20[3] ^ sign), global_second} : {(in_data_20[3] ^ sign), global_min};
        out_data_21 = (in_data_21[2:0] == global_min) ? {(in_data_21[3] ^ sign), global_second} : {(in_data_21[3] ^ sign), global_min};
        out_data_22 = (in_data_22[2:0] == global_min) ? {(in_data_22[3] ^ sign), global_second} : {(in_data_22[3] ^ sign), global_min};
        out_data_23 = (in_data_23[2:0] == global_min) ? {(in_data_23[3] ^ sign), global_second} : {(in_data_23[3] ^ sign), global_min};
        out_data_24 = (in_data_24[2:0] == global_min) ? {(in_data_24[3] ^ sign), global_second} : {(in_data_24[3] ^ sign), global_min};
        out_data_25 = (in_data_25[2:0] == global_min) ? {(in_data_25[3] ^ sign), global_second} : {(in_data_25[3] ^ sign), global_min};
        out_data_26 = (in_data_26[2:0] == global_min) ? {(in_data_26[3] ^ sign), global_second} : {(in_data_26[3] ^ sign), global_min};
        out_data_27 = (in_data_27[2:0] == global_min) ? {(in_data_27[3] ^ sign), global_second} : {(in_data_27[3] ^ sign), global_min};
        out_data_28 = (in_data_28[2:0] == global_min) ? {(in_data_28[3] ^ sign), global_second} : {(in_data_28[3] ^ sign), global_min};
        out_data_29 = (in_data_29[2:0] == global_min) ? {(in_data_29[3] ^ sign), global_second} : {(in_data_29[3] ^ sign), global_min};
        out_data_30 = (in_data_30[2:0] == global_min) ? {(in_data_30[3] ^ sign), global_second} : {(in_data_30[3] ^ sign), global_min};
        out_data_31 = (in_data_31[2:0] == global_min) ? {(in_data_31[3] ^ sign), global_second} : {(in_data_31[3] ^ sign), global_min};
        out_data_32 = (in_data_32[2:0] == global_min) ? {(in_data_32[3] ^ sign), global_second} : {(in_data_32[3] ^ sign), global_min};
        out_data_33 = (in_data_33[2:0] == global_min) ? {(in_data_33[3] ^ sign), global_second} : {(in_data_33[3] ^ sign), global_min};
        out_data_34 = (in_data_34[2:0] == global_min) ? {(in_data_34[3] ^ sign), global_second} : {(in_data_34[3] ^ sign), global_min};
        out_data_35 = (in_data_35[2:0] == global_min) ? {(in_data_35[3] ^ sign), global_second} : {(in_data_35[3] ^ sign), global_min};
        out_data_36 = (in_data_36[2:0] == global_min) ? {(in_data_36[3] ^ sign), global_second} : {(in_data_36[3] ^ sign), global_min};
        out_data_37 = (in_data_37[2:0] == global_min) ? {(in_data_37[3] ^ sign), global_second} : {(in_data_37[3] ^ sign), global_min};
        out_data_38 = (in_data_38[2:0] == global_min) ? {(in_data_38[3] ^ sign), global_second} : {(in_data_38[3] ^ sign), global_min};
        out_data_39 = (in_data_39[2:0] == global_min) ? {(in_data_39[3] ^ sign), global_second} : {(in_data_39[3] ^ sign), global_min};
        out_data_40 = (in_data_40[2:0] == global_min) ? {(in_data_40[3] ^ sign), global_second} : {(in_data_40[3] ^ sign), global_min};
        out_data_41 = (in_data_41[2:0] == global_min) ? {(in_data_41[3] ^ sign), global_second} : {(in_data_41[3] ^ sign), global_min};
        out_data_42 = (in_data_42[2:0] == global_min) ? {(in_data_42[3] ^ sign), global_second} : {(in_data_42[3] ^ sign), global_min};
        out_data_43 = (in_data_43[2:0] == global_min) ? {(in_data_43[3] ^ sign), global_second} : {(in_data_43[3] ^ sign), global_min};
        out_data_44 = (in_data_44[2:0] == global_min) ? {(in_data_44[3] ^ sign), global_second} : {(in_data_44[3] ^ sign), global_min};
        out_data_45 = (in_data_45[2:0] == global_min) ? {(in_data_45[3] ^ sign), global_second} : {(in_data_45[3] ^ sign), global_min};
        out_data_46 = (in_data_46[2:0] == global_min) ? {(in_data_46[3] ^ sign), global_second} : {(in_data_46[3] ^ sign), global_min};
        out_data_47 = (in_data_47[2:0] == global_min) ? {(in_data_47[3] ^ sign), global_second} : {(in_data_47[3] ^ sign), global_min};
        out_data_48 = (in_data_48[2:0] == global_min) ? {(in_data_48[3] ^ sign), global_second} : {(in_data_48[3] ^ sign), global_min};
        out_data_49 = (in_data_49[2:0] == global_min) ? {(in_data_49[3] ^ sign), global_second} : {(in_data_49[3] ^ sign), global_min};
        out_data_50 = (in_data_50[2:0] == global_min) ? {(in_data_50[3] ^ sign), global_second} : {(in_data_50[3] ^ sign), global_min};
        out_data_51 = (in_data_51[2:0] == global_min) ? {(in_data_51[3] ^ sign), global_second} : {(in_data_51[3] ^ sign), global_min};
        out_data_52 = (in_data_52[2:0] == global_min) ? {(in_data_52[3] ^ sign), global_second} : {(in_data_52[3] ^ sign), global_min};
        out_data_53 = (in_data_53[2:0] == global_min) ? {(in_data_53[3] ^ sign), global_second} : {(in_data_53[3] ^ sign), global_min};
        out_data_54 = (in_data_54[2:0] == global_min) ? {(in_data_54[3] ^ sign), global_second} : {(in_data_54[3] ^ sign), global_min};
        out_data_55 = (in_data_55[2:0] == global_min) ? {(in_data_55[3] ^ sign), global_second} : {(in_data_55[3] ^ sign), global_min};
        out_data_56 = (in_data_56[2:0] == global_min) ? {(in_data_56[3] ^ sign), global_second} : {(in_data_56[3] ^ sign), global_min};
        out_data_57 = (in_data_57[2:0] == global_min) ? {(in_data_57[3] ^ sign), global_second} : {(in_data_57[3] ^ sign), global_min};
        out_data_58 = (in_data_58[2:0] == global_min) ? {(in_data_58[3] ^ sign), global_second} : {(in_data_58[3] ^ sign), global_min};
        out_data_59 = (in_data_59[2:0] == global_min) ? {(in_data_59[3] ^ sign), global_second} : {(in_data_59[3] ^ sign), global_min};
        out_data_60 = (in_data_60[2:0] == global_min) ? {(in_data_60[3] ^ sign), global_second} : {(in_data_60[3] ^ sign), global_min};
        out_data_61 = (in_data_61[2:0] == global_min) ? {(in_data_61[3] ^ sign), global_second} : {(in_data_61[3] ^ sign), global_min};
        out_data_62 = (in_data_62[2:0] == global_min) ? {(in_data_62[3] ^ sign), global_second} : {(in_data_62[3] ^ sign), global_min};
        out_data_63 = (in_data_63[2:0] == global_min) ? {(in_data_63[3] ^ sign), global_second} : {(in_data_63[3] ^ sign), global_min};
        out_data_64 = (in_data_64[2:0] == global_min) ? {(in_data_64[3] ^ sign), global_second} : {(in_data_64[3] ^ sign), global_min};
        out_data_65 = (in_data_65[2:0] == global_min) ? {(in_data_65[3] ^ sign), global_second} : {(in_data_65[3] ^ sign), global_min};
        out_data_66 = (in_data_66[2:0] == global_min) ? {(in_data_66[3] ^ sign), global_second} : {(in_data_66[3] ^ sign), global_min};
        out_data_67 = (in_data_67[2:0] == global_min) ? {(in_data_67[3] ^ sign), global_second} : {(in_data_67[3] ^ sign), global_min};
        out_data_68 = (in_data_68[2:0] == global_min) ? {(in_data_68[3] ^ sign), global_second} : {(in_data_68[3] ^ sign), global_min};
        out_data_69 = (in_data_69[2:0] == global_min) ? {(in_data_69[3] ^ sign), global_second} : {(in_data_69[3] ^ sign), global_min};
        out_data_70 = (in_data_70[2:0] == global_min) ? {(in_data_70[3] ^ sign), global_second} : {(in_data_70[3] ^ sign), global_min};
        out_data_71 = (in_data_71[2:0] == global_min) ? {(in_data_71[3] ^ sign), global_second} : {(in_data_71[3] ^ sign), global_min};
        out_data_72 = (in_data_72[2:0] == global_min) ? {(in_data_72[3] ^ sign), global_second} : {(in_data_72[3] ^ sign), global_min};
        out_data_73 = (in_data_73[2:0] == global_min) ? {(in_data_73[3] ^ sign), global_second} : {(in_data_73[3] ^ sign), global_min};
        out_data_74 = (in_data_74[2:0] == global_min) ? {(in_data_74[3] ^ sign), global_second} : {(in_data_74[3] ^ sign), global_min};
        out_data_75 = (in_data_75[2:0] == global_min) ? {(in_data_75[3] ^ sign), global_second} : {(in_data_75[3] ^ sign), global_min};
        out_data_76 = (in_data_76[2:0] == global_min) ? {(in_data_76[3] ^ sign), global_second} : {(in_data_76[3] ^ sign), global_min};
        out_data_77 = (in_data_77[2:0] == global_min) ? {(in_data_77[3] ^ sign), global_second} : {(in_data_77[3] ^ sign), global_min};
        out_data_78 = (in_data_78[2:0] == global_min) ? {(in_data_78[3] ^ sign), global_second} : {(in_data_78[3] ^ sign), global_min};
        out_data_79 = (in_data_79[2:0] == global_min) ? {(in_data_79[3] ^ sign), global_second} : {(in_data_79[3] ^ sign), global_min};
        out_data_80 = (in_data_80[2:0] == global_min) ? {(in_data_80[3] ^ sign), global_second} : {(in_data_80[3] ^ sign), global_min};
        out_data_81 = (in_data_81[2:0] == global_min) ? {(in_data_81[3] ^ sign), global_second} : {(in_data_81[3] ^ sign), global_min};
        out_data_82 = (in_data_82[2:0] == global_min) ? {(in_data_82[3] ^ sign), global_second} : {(in_data_82[3] ^ sign), global_min};
        out_data_83 = (in_data_83[2:0] == global_min) ? {(in_data_83[3] ^ sign), global_second} : {(in_data_83[3] ^ sign), global_min};
        out_data_84 = (in_data_84[2:0] == global_min) ? {(in_data_84[3] ^ sign), global_second} : {(in_data_84[3] ^ sign), global_min};
        out_data_85 = (in_data_85[2:0] == global_min) ? {(in_data_85[3] ^ sign), global_second} : {(in_data_85[3] ^ sign), global_min};
        out_data_86 = (in_data_86[2:0] == global_min) ? {(in_data_86[3] ^ sign), global_second} : {(in_data_86[3] ^ sign), global_min};
        out_data_87 = (in_data_87[2:0] == global_min) ? {(in_data_87[3] ^ sign), global_second} : {(in_data_87[3] ^ sign), global_min};
        out_data_88 = (in_data_88[2:0] == global_min) ? {(in_data_88[3] ^ sign), global_second} : {(in_data_88[3] ^ sign), global_min};
        out_data_89 = (in_data_89[2:0] == global_min) ? {(in_data_89[3] ^ sign), global_second} : {(in_data_89[3] ^ sign), global_min};
        out_data_90 = (in_data_90[2:0] == global_min) ? {(in_data_90[3] ^ sign), global_second} : {(in_data_90[3] ^ sign), global_min};
        out_data_91 = (in_data_91[2:0] == global_min) ? {(in_data_91[3] ^ sign), global_second} : {(in_data_91[3] ^ sign), global_min};
        out_data_92 = (in_data_92[2:0] == global_min) ? {(in_data_92[3] ^ sign), global_second} : {(in_data_92[3] ^ sign), global_min};
        out_data_93 = (in_data_93[2:0] == global_min) ? {(in_data_93[3] ^ sign), global_second} : {(in_data_93[3] ^ sign), global_min};
        out_data_94 = (in_data_94[2:0] == global_min) ? {(in_data_94[3] ^ sign), global_second} : {(in_data_94[3] ^ sign), global_min};
        out_data_95 = (in_data_95[2:0] == global_min) ? {(in_data_95[3] ^ sign), global_second} : {(in_data_95[3] ^ sign), global_min};
        out_data_96 = (in_data_96[2:0] == global_min) ? {(in_data_96[3] ^ sign), global_second} : {(in_data_96[3] ^ sign), global_min};
        out_data_97 = (in_data_97[2:0] == global_min) ? {(in_data_97[3] ^ sign), global_second} : {(in_data_97[3] ^ sign), global_min};
        out_data_98 = (in_data_98[2:0] == global_min) ? {(in_data_98[3] ^ sign), global_second} : {(in_data_98[3] ^ sign), global_min};
        out_data_99 = (in_data_99[2:0] == global_min) ? {(in_data_99[3] ^ sign), global_second} : {(in_data_99[3] ^ sign), global_min};
        out_data_100 = (in_data_100[2:0] == global_min) ? {(in_data_100[3] ^ sign), global_second} : {(in_data_100[3] ^ sign), global_min};
        out_data_101 = (in_data_101[2:0] == global_min) ? {(in_data_101[3] ^ sign), global_second} : {(in_data_101[3] ^ sign), global_min};
        out_data_102 = (in_data_102[2:0] == global_min) ? {(in_data_102[3] ^ sign), global_second} : {(in_data_102[3] ^ sign), global_min};
    end

endmodule