module buffer_in #(
        parameter QNT_BIT            = 4,  // LLR量化位宽为4位
        parameter QC_LDPC_COL_COUNT  = 533,  // 基矩阵列数
    parameter QC_LDPC_BLOCK_SIZE = 64   // 扩展因子
    ) (
        input wire               sys_clk,
        input wire               sys_rst_n,
        input wire               sink_star,          // 输入开始
        input wire               sink_stop,          // 输入停止
        input wire [QNT_BIT-1:0] sink,               // 输入数据
        input wire               flag_org_update,    // 写入下一帧

        output reg                buffer_wr_en,     // 给后面 combine_ram_llr 的写入 en 信号
        output wire [QNT_BIT-1:0] rr_data_1,       // 读取数据
        output wire [QNT_BIT-1:0] rr_data_2,
        output wire [QNT_BIT-1:0] rr_data_3,
        output wire [QNT_BIT-1:0] rr_data_4,
        output wire [QNT_BIT-1:0] rr_data_5,
        output wire [QNT_BIT-1:0] rr_data_6,
        output wire [QNT_BIT-1:0] rr_data_7,
        output wire [QNT_BIT-1:0] rr_data_8,
        output wire [QNT_BIT-1:0] rr_data_9,
        output wire [QNT_BIT-1:0] rr_data_10,
        output wire [QNT_BIT-1:0] rr_data_11,
        output wire [QNT_BIT-1:0] rr_data_12,
        output wire [QNT_BIT-1:0] rr_data_13,
        output wire [QNT_BIT-1:0] rr_data_14,
        output wire [QNT_BIT-1:0] rr_data_15,
        output wire [QNT_BIT-1:0] rr_data_16,
        output wire [QNT_BIT-1:0] rr_data_17,
        output wire [QNT_BIT-1:0] rr_data_18,
        output wire [QNT_BIT-1:0] rr_data_19,
        output wire [QNT_BIT-1:0] rr_data_20,
        output wire [QNT_BIT-1:0] rr_data_21,
        output wire [QNT_BIT-1:0] rr_data_22,
        output wire [QNT_BIT-1:0] rr_data_23,
        output wire [QNT_BIT-1:0] rr_data_24,
        output wire [QNT_BIT-1:0] rr_data_25,
        output wire [QNT_BIT-1:0] rr_data_26,
        output wire [QNT_BIT-1:0] rr_data_27,
        output wire [QNT_BIT-1:0] rr_data_28,
        output wire [QNT_BIT-1:0] rr_data_29,
        output wire [QNT_BIT-1:0] rr_data_30,
        output wire [QNT_BIT-1:0] rr_data_31,
        output wire [QNT_BIT-1:0] rr_data_32,
        output wire [QNT_BIT-1:0] rr_data_33,
        output wire [QNT_BIT-1:0] rr_data_34,
        output wire [QNT_BIT-1:0] rr_data_35,
        output wire [QNT_BIT-1:0] rr_data_36,
        output wire [QNT_BIT-1:0] rr_data_37,
        output wire [QNT_BIT-1:0] rr_data_38,
        output wire [QNT_BIT-1:0] rr_data_39,
        output wire [QNT_BIT-1:0] rr_data_40,
        output wire [QNT_BIT-1:0] rr_data_41,
        output wire [QNT_BIT-1:0] rr_data_42,
        output wire [QNT_BIT-1:0] rr_data_43,
        output wire [QNT_BIT-1:0] rr_data_44,
        output wire [QNT_BIT-1:0] rr_data_45,
        output wire [QNT_BIT-1:0] rr_data_46,
        output wire [QNT_BIT-1:0] rr_data_47,
        output wire [QNT_BIT-1:0] rr_data_48,
        output wire [QNT_BIT-1:0] rr_data_49,
        output wire [QNT_BIT-1:0] rr_data_50,
        output wire [QNT_BIT-1:0] rr_data_51,
        output wire [QNT_BIT-1:0] rr_data_52,
        output wire [QNT_BIT-1:0] rr_data_53,
        output wire [QNT_BIT-1:0] rr_data_54,
        output wire [QNT_BIT-1:0] rr_data_55,
        output wire [QNT_BIT-1:0] rr_data_56,
        output wire [QNT_BIT-1:0] rr_data_57,
        output wire [QNT_BIT-1:0] rr_data_58,
        output wire [QNT_BIT-1:0] rr_data_59,
        output wire [QNT_BIT-1:0] rr_data_60,
        output wire [QNT_BIT-1:0] rr_data_61,
        output wire [QNT_BIT-1:0] rr_data_62,
        output wire [QNT_BIT-1:0] rr_data_63,
        output wire [QNT_BIT-1:0] rr_data_64,
        output wire [QNT_BIT-1:0] rr_data_65,
        output wire [QNT_BIT-1:0] rr_data_66,
        output wire [QNT_BIT-1:0] rr_data_67,
        output wire [QNT_BIT-1:0] rr_data_68,
        output wire [QNT_BIT-1:0] rr_data_69,
        output wire [QNT_BIT-1:0] rr_data_70,
        output wire [QNT_BIT-1:0] rr_data_71,
        output wire [QNT_BIT-1:0] rr_data_72,
        output wire [QNT_BIT-1:0] rr_data_73,
        output wire [QNT_BIT-1:0] rr_data_74,
        output wire [QNT_BIT-1:0] rr_data_75,
        output wire [QNT_BIT-1:0] rr_data_76,
        output wire [QNT_BIT-1:0] rr_data_77,
        output wire [QNT_BIT-1:0] rr_data_78,
        output wire [QNT_BIT-1:0] rr_data_79,
        output wire [QNT_BIT-1:0] rr_data_80,
        output wire [QNT_BIT-1:0] rr_data_81,
        output wire [QNT_BIT-1:0] rr_data_82,
        output wire [QNT_BIT-1:0] rr_data_83,
        output wire [QNT_BIT-1:0] rr_data_84,
        output wire [QNT_BIT-1:0] rr_data_85,
        output wire [QNT_BIT-1:0] rr_data_86,
        output wire [QNT_BIT-1:0] rr_data_87,
        output wire [QNT_BIT-1:0] rr_data_88,
        output wire [QNT_BIT-1:0] rr_data_89,
        output wire [QNT_BIT-1:0] rr_data_90,
        output wire [QNT_BIT-1:0] rr_data_91,
        output wire [QNT_BIT-1:0] rr_data_92,
        output wire [QNT_BIT-1:0] rr_data_93,
        output wire [QNT_BIT-1:0] rr_data_94,
        output wire [QNT_BIT-1:0] rr_data_95,
        output wire [QNT_BIT-1:0] rr_data_96,
        output wire [QNT_BIT-1:0] rr_data_97,
        output wire [QNT_BIT-1:0] rr_data_98,
        output wire [QNT_BIT-1:0] rr_data_99,
        output wire [QNT_BIT-1:0] rr_data_100,
        output wire [QNT_BIT-1:0] rr_data_101,
        output wire [QNT_BIT-1:0] rr_data_102,
        output wire [QNT_BIT-1:0] rr_data_103,
        output wire [QNT_BIT-1:0] rr_data_104,
        output wire [QNT_BIT-1:0] rr_data_105,
        output wire [QNT_BIT-1:0] rr_data_106,
        output wire [QNT_BIT-1:0] rr_data_107,
        output wire [QNT_BIT-1:0] rr_data_108,
        output wire [QNT_BIT-1:0] rr_data_109,
        output wire [QNT_BIT-1:0] rr_data_110,
        output wire [QNT_BIT-1:0] rr_data_111,
        output wire [QNT_BIT-1:0] rr_data_112,
        output wire [QNT_BIT-1:0] rr_data_113,
        output wire [QNT_BIT-1:0] rr_data_114,
        output wire [QNT_BIT-1:0] rr_data_115,
        output wire [QNT_BIT-1:0] rr_data_116,
        output wire [QNT_BIT-1:0] rr_data_117,
        output wire [QNT_BIT-1:0] rr_data_118,
        output wire [QNT_BIT-1:0] rr_data_119,
        output wire [QNT_BIT-1:0] rr_data_120,
        output wire [QNT_BIT-1:0] rr_data_121,
        output wire [QNT_BIT-1:0] rr_data_122,
        output wire [QNT_BIT-1:0] rr_data_123,
        output wire [QNT_BIT-1:0] rr_data_124,
        output wire [QNT_BIT-1:0] rr_data_125,
        output wire [QNT_BIT-1:0] rr_data_126,
        output wire [QNT_BIT-1:0] rr_data_127,
        output wire [QNT_BIT-1:0] rr_data_128,
        output wire [QNT_BIT-1:0] rr_data_129,
        output wire [QNT_BIT-1:0] rr_data_130,
        output wire [QNT_BIT-1:0] rr_data_131,
        output wire [QNT_BIT-1:0] rr_data_132,
        output wire [QNT_BIT-1:0] rr_data_133,
        output wire [QNT_BIT-1:0] rr_data_134,
        output wire [QNT_BIT-1:0] rr_data_135,
        output wire [QNT_BIT-1:0] rr_data_136,
        output wire [QNT_BIT-1:0] rr_data_137,
        output wire [QNT_BIT-1:0] rr_data_138,
        output wire [QNT_BIT-1:0] rr_data_139,
        output wire [QNT_BIT-1:0] rr_data_140,
        output wire [QNT_BIT-1:0] rr_data_141,
        output wire [QNT_BIT-1:0] rr_data_142,
        output wire [QNT_BIT-1:0] rr_data_143,
        output wire [QNT_BIT-1:0] rr_data_144,
        output wire [QNT_BIT-1:0] rr_data_145,
        output wire [QNT_BIT-1:0] rr_data_146,
        output wire [QNT_BIT-1:0] rr_data_147,
        output wire [QNT_BIT-1:0] rr_data_148,
        output wire [QNT_BIT-1:0] rr_data_149,
        output wire [QNT_BIT-1:0] rr_data_150,
        output wire [QNT_BIT-1:0] rr_data_151,
        output wire [QNT_BIT-1:0] rr_data_152,
        output wire [QNT_BIT-1:0] rr_data_153,
        output wire [QNT_BIT-1:0] rr_data_154,
        output wire [QNT_BIT-1:0] rr_data_155,
        output wire [QNT_BIT-1:0] rr_data_156,
        output wire [QNT_BIT-1:0] rr_data_157,
        output wire [QNT_BIT-1:0] rr_data_158,
        output wire [QNT_BIT-1:0] rr_data_159,
        output wire [QNT_BIT-1:0] rr_data_160,
        output wire [QNT_BIT-1:0] rr_data_161,
        output wire [QNT_BIT-1:0] rr_data_162,
        output wire [QNT_BIT-1:0] rr_data_163,
        output wire [QNT_BIT-1:0] rr_data_164,
        output wire [QNT_BIT-1:0] rr_data_165,
        output wire [QNT_BIT-1:0] rr_data_166,
        output wire [QNT_BIT-1:0] rr_data_167,
        output wire [QNT_BIT-1:0] rr_data_168,
        output wire [QNT_BIT-1:0] rr_data_169,
        output wire [QNT_BIT-1:0] rr_data_170,
        output wire [QNT_BIT-1:0] rr_data_171,
        output wire [QNT_BIT-1:0] rr_data_172,
        output wire [QNT_BIT-1:0] rr_data_173,
        output wire [QNT_BIT-1:0] rr_data_174,
        output wire [QNT_BIT-1:0] rr_data_175,
        output wire [QNT_BIT-1:0] rr_data_176,
        output wire [QNT_BIT-1:0] rr_data_177,
        output wire [QNT_BIT-1:0] rr_data_178,
        output wire [QNT_BIT-1:0] rr_data_179,
        output wire [QNT_BIT-1:0] rr_data_180,
        output wire [QNT_BIT-1:0] rr_data_181,
        output wire [QNT_BIT-1:0] rr_data_182,
        output wire [QNT_BIT-1:0] rr_data_183,
        output wire [QNT_BIT-1:0] rr_data_184,
        output wire [QNT_BIT-1:0] rr_data_185,
        output wire [QNT_BIT-1:0] rr_data_186,
        output wire [QNT_BIT-1:0] rr_data_187,
        output wire [QNT_BIT-1:0] rr_data_188,
        output wire [QNT_BIT-1:0] rr_data_189,
        output wire [QNT_BIT-1:0] rr_data_190,
        output wire [QNT_BIT-1:0] rr_data_191,
        output wire [QNT_BIT-1:0] rr_data_192,
        output wire [QNT_BIT-1:0] rr_data_193,
        output wire [QNT_BIT-1:0] rr_data_194,
        output wire [QNT_BIT-1:0] rr_data_195,
        output wire [QNT_BIT-1:0] rr_data_196,
        output wire [QNT_BIT-1:0] rr_data_197,
        output wire [QNT_BIT-1:0] rr_data_198,
        output wire [QNT_BIT-1:0] rr_data_199,
        output wire [QNT_BIT-1:0] rr_data_200,
        output wire [QNT_BIT-1:0] rr_data_201,
        output wire [QNT_BIT-1:0] rr_data_202,
        output wire [QNT_BIT-1:0] rr_data_203,
        output wire [QNT_BIT-1:0] rr_data_204,
        output wire [QNT_BIT-1:0] rr_data_205,
        output wire [QNT_BIT-1:0] rr_data_206,
        output wire [QNT_BIT-1:0] rr_data_207,
        output wire [QNT_BIT-1:0] rr_data_208,
        output wire [QNT_BIT-1:0] rr_data_209,
        output wire [QNT_BIT-1:0] rr_data_210,
        output wire [QNT_BIT-1:0] rr_data_211,
        output wire [QNT_BIT-1:0] rr_data_212,
        output wire [QNT_BIT-1:0] rr_data_213,
        output wire [QNT_BIT-1:0] rr_data_214,
        output wire [QNT_BIT-1:0] rr_data_215,
        output wire [QNT_BIT-1:0] rr_data_216,
        output wire [QNT_BIT-1:0] rr_data_217,
        output wire [QNT_BIT-1:0] rr_data_218,
        output wire [QNT_BIT-1:0] rr_data_219,
        output wire [QNT_BIT-1:0] rr_data_220,
        output wire [QNT_BIT-1:0] rr_data_221,
        output wire [QNT_BIT-1:0] rr_data_222,
        output wire [QNT_BIT-1:0] rr_data_223,
        output wire [QNT_BIT-1:0] rr_data_224,
        output wire [QNT_BIT-1:0] rr_data_225,
        output wire [QNT_BIT-1:0] rr_data_226,
        output wire [QNT_BIT-1:0] rr_data_227,
        output wire [QNT_BIT-1:0] rr_data_228,
        output wire [QNT_BIT-1:0] rr_data_229,
        output wire [QNT_BIT-1:0] rr_data_230,
        output wire [QNT_BIT-1:0] rr_data_231,
        output wire [QNT_BIT-1:0] rr_data_232,
        output wire [QNT_BIT-1:0] rr_data_233,
        output wire [QNT_BIT-1:0] rr_data_234,
        output wire [QNT_BIT-1:0] rr_data_235,
        output wire [QNT_BIT-1:0] rr_data_236,
        output wire [QNT_BIT-1:0] rr_data_237,
        output wire [QNT_BIT-1:0] rr_data_238,
        output wire [QNT_BIT-1:0] rr_data_239,
        output wire [QNT_BIT-1:0] rr_data_240,
        output wire [QNT_BIT-1:0] rr_data_241,
        output wire [QNT_BIT-1:0] rr_data_242,
        output wire [QNT_BIT-1:0] rr_data_243,
        output wire [QNT_BIT-1:0] rr_data_244,
        output wire [QNT_BIT-1:0] rr_data_245,
        output wire [QNT_BIT-1:0] rr_data_246,
        output wire [QNT_BIT-1:0] rr_data_247,
        output wire [QNT_BIT-1:0] rr_data_248,
        output wire [QNT_BIT-1:0] rr_data_249,
        output wire [QNT_BIT-1:0] rr_data_250,
        output wire [QNT_BIT-1:0] rr_data_251,
        output wire [QNT_BIT-1:0] rr_data_252,
        output wire [QNT_BIT-1:0] rr_data_253,
        output wire [QNT_BIT-1:0] rr_data_254,
        output wire [QNT_BIT-1:0] rr_data_255,
        output wire [QNT_BIT-1:0] rr_data_256,
        output wire [QNT_BIT-1:0] rr_data_257,
        output wire [QNT_BIT-1:0] rr_data_258,
        output wire [QNT_BIT-1:0] rr_data_259,
        output wire [QNT_BIT-1:0] rr_data_260,
        output wire [QNT_BIT-1:0] rr_data_261,
        output wire [QNT_BIT-1:0] rr_data_262,
        output wire [QNT_BIT-1:0] rr_data_263,
        output wire [QNT_BIT-1:0] rr_data_264,
        output wire [QNT_BIT-1:0] rr_data_265,
        output wire [QNT_BIT-1:0] rr_data_266,
        output wire [QNT_BIT-1:0] rr_data_267,
        output wire [QNT_BIT-1:0] rr_data_268,
        output wire [QNT_BIT-1:0] rr_data_269,
        output wire [QNT_BIT-1:0] rr_data_270,
        output wire [QNT_BIT-1:0] rr_data_271,
        output wire [QNT_BIT-1:0] rr_data_272,
        output wire [QNT_BIT-1:0] rr_data_273,
        output wire [QNT_BIT-1:0] rr_data_274,
        output wire [QNT_BIT-1:0] rr_data_275,
        output wire [QNT_BIT-1:0] rr_data_276,
        output wire [QNT_BIT-1:0] rr_data_277,
        output wire [QNT_BIT-1:0] rr_data_278,
        output wire [QNT_BIT-1:0] rr_data_279,
        output wire [QNT_BIT-1:0] rr_data_280,
        output wire [QNT_BIT-1:0] rr_data_281,
        output wire [QNT_BIT-1:0] rr_data_282,
        output wire [QNT_BIT-1:0] rr_data_283,
        output wire [QNT_BIT-1:0] rr_data_284,
        output wire [QNT_BIT-1:0] rr_data_285,
        output wire [QNT_BIT-1:0] rr_data_286,
        output wire [QNT_BIT-1:0] rr_data_287,
        output wire [QNT_BIT-1:0] rr_data_288,
        output wire [QNT_BIT-1:0] rr_data_289,
        output wire [QNT_BIT-1:0] rr_data_290,
        output wire [QNT_BIT-1:0] rr_data_291,
        output wire [QNT_BIT-1:0] rr_data_292,
        output wire [QNT_BIT-1:0] rr_data_293,
        output wire [QNT_BIT-1:0] rr_data_294,
        output wire [QNT_BIT-1:0] rr_data_295,
        output wire [QNT_BIT-1:0] rr_data_296,
        output wire [QNT_BIT-1:0] rr_data_297,
        output wire [QNT_BIT-1:0] rr_data_298,
        output wire [QNT_BIT-1:0] rr_data_299,
        output wire [QNT_BIT-1:0] rr_data_300,
        output wire [QNT_BIT-1:0] rr_data_301,
        output wire [QNT_BIT-1:0] rr_data_302,
        output wire [QNT_BIT-1:0] rr_data_303,
        output wire [QNT_BIT-1:0] rr_data_304,
        output wire [QNT_BIT-1:0] rr_data_305,
        output wire [QNT_BIT-1:0] rr_data_306,
        output wire [QNT_BIT-1:0] rr_data_307,
        output wire [QNT_BIT-1:0] rr_data_308,
        output wire [QNT_BIT-1:0] rr_data_309,
        output wire [QNT_BIT-1:0] rr_data_310,
        output wire [QNT_BIT-1:0] rr_data_311,
        output wire [QNT_BIT-1:0] rr_data_312,
        output wire [QNT_BIT-1:0] rr_data_313,
        output wire [QNT_BIT-1:0] rr_data_314,
        output wire [QNT_BIT-1:0] rr_data_315,
        output wire [QNT_BIT-1:0] rr_data_316,
        output wire [QNT_BIT-1:0] rr_data_317,
        output wire [QNT_BIT-1:0] rr_data_318,
        output wire [QNT_BIT-1:0] rr_data_319,
        output wire [QNT_BIT-1:0] rr_data_320,
        output wire [QNT_BIT-1:0] rr_data_321,
        output wire [QNT_BIT-1:0] rr_data_322,
        output wire [QNT_BIT-1:0] rr_data_323,
        output wire [QNT_BIT-1:0] rr_data_324,
        output wire [QNT_BIT-1:0] rr_data_325,
        output wire [QNT_BIT-1:0] rr_data_326,
        output wire [QNT_BIT-1:0] rr_data_327,
        output wire [QNT_BIT-1:0] rr_data_328,
        output wire [QNT_BIT-1:0] rr_data_329,
        output wire [QNT_BIT-1:0] rr_data_330,
        output wire [QNT_BIT-1:0] rr_data_331,
        output wire [QNT_BIT-1:0] rr_data_332,
        output wire [QNT_BIT-1:0] rr_data_333,
        output wire [QNT_BIT-1:0] rr_data_334,
        output wire [QNT_BIT-1:0] rr_data_335,
        output wire [QNT_BIT-1:0] rr_data_336,
        output wire [QNT_BIT-1:0] rr_data_337,
        output wire [QNT_BIT-1:0] rr_data_338,
        output wire [QNT_BIT-1:0] rr_data_339,
        output wire [QNT_BIT-1:0] rr_data_340,
        output wire [QNT_BIT-1:0] rr_data_341,
        output wire [QNT_BIT-1:0] rr_data_342,
        output wire [QNT_BIT-1:0] rr_data_343,
        output wire [QNT_BIT-1:0] rr_data_344,
        output wire [QNT_BIT-1:0] rr_data_345,
        output wire [QNT_BIT-1:0] rr_data_346,
        output wire [QNT_BIT-1:0] rr_data_347,
        output wire [QNT_BIT-1:0] rr_data_348,
        output wire [QNT_BIT-1:0] rr_data_349,
        output wire [QNT_BIT-1:0] rr_data_350,
        output wire [QNT_BIT-1:0] rr_data_351,
        output wire [QNT_BIT-1:0] rr_data_352,
        output wire [QNT_BIT-1:0] rr_data_353,
        output wire [QNT_BIT-1:0] rr_data_354,
        output wire [QNT_BIT-1:0] rr_data_355,
        output wire [QNT_BIT-1:0] rr_data_356,
        output wire [QNT_BIT-1:0] rr_data_357,
        output wire [QNT_BIT-1:0] rr_data_358,
        output wire [QNT_BIT-1:0] rr_data_359,
        output wire [QNT_BIT-1:0] rr_data_360,
        output wire [QNT_BIT-1:0] rr_data_361,
        output wire [QNT_BIT-1:0] rr_data_362,
        output wire [QNT_BIT-1:0] rr_data_363,
        output wire [QNT_BIT-1:0] rr_data_364,
        output wire [QNT_BIT-1:0] rr_data_365,
        output wire [QNT_BIT-1:0] rr_data_366,
        output wire [QNT_BIT-1:0] rr_data_367,
        output wire [QNT_BIT-1:0] rr_data_368,
        output wire [QNT_BIT-1:0] rr_data_369,
        output wire [QNT_BIT-1:0] rr_data_370,
        output wire [QNT_BIT-1:0] rr_data_371,
        output wire [QNT_BIT-1:0] rr_data_372,
        output wire [QNT_BIT-1:0] rr_data_373,
        output wire [QNT_BIT-1:0] rr_data_374,
        output wire [QNT_BIT-1:0] rr_data_375,
        output wire [QNT_BIT-1:0] rr_data_376,
        output wire [QNT_BIT-1:0] rr_data_377,
        output wire [QNT_BIT-1:0] rr_data_378,
        output wire [QNT_BIT-1:0] rr_data_379,
        output wire [QNT_BIT-1:0] rr_data_380,
        output wire [QNT_BIT-1:0] rr_data_381,
        output wire [QNT_BIT-1:0] rr_data_382,
        output wire [QNT_BIT-1:0] rr_data_383,
        output wire [QNT_BIT-1:0] rr_data_384,
        output wire [QNT_BIT-1:0] rr_data_385,
        output wire [QNT_BIT-1:0] rr_data_386,
        output wire [QNT_BIT-1:0] rr_data_387,
        output wire [QNT_BIT-1:0] rr_data_388,
        output wire [QNT_BIT-1:0] rr_data_389,
        output wire [QNT_BIT-1:0] rr_data_390,
        output wire [QNT_BIT-1:0] rr_data_391,
        output wire [QNT_BIT-1:0] rr_data_392,
        output wire [QNT_BIT-1:0] rr_data_393,
        output wire [QNT_BIT-1:0] rr_data_394,
        output wire [QNT_BIT-1:0] rr_data_395,
        output wire [QNT_BIT-1:0] rr_data_396,
        output wire [QNT_BIT-1:0] rr_data_397,
        output wire [QNT_BIT-1:0] rr_data_398,
        output wire [QNT_BIT-1:0] rr_data_399,
        output wire [QNT_BIT-1:0] rr_data_400,
        output wire [QNT_BIT-1:0] rr_data_401,
        output wire [QNT_BIT-1:0] rr_data_402,
        output wire [QNT_BIT-1:0] rr_data_403,
        output wire [QNT_BIT-1:0] rr_data_404,
        output wire [QNT_BIT-1:0] rr_data_405,
        output wire [QNT_BIT-1:0] rr_data_406,
        output wire [QNT_BIT-1:0] rr_data_407,
        output wire [QNT_BIT-1:0] rr_data_408,
        output wire [QNT_BIT-1:0] rr_data_409,
        output wire [QNT_BIT-1:0] rr_data_410,
        output wire [QNT_BIT-1:0] rr_data_411,
        output wire [QNT_BIT-1:0] rr_data_412,
        output wire [QNT_BIT-1:0] rr_data_413,
        output wire [QNT_BIT-1:0] rr_data_414,
        output wire [QNT_BIT-1:0] rr_data_415,
        output wire [QNT_BIT-1:0] rr_data_416,
        output wire [QNT_BIT-1:0] rr_data_417,
        output wire [QNT_BIT-1:0] rr_data_418,
        output wire [QNT_BIT-1:0] rr_data_419,
        output wire [QNT_BIT-1:0] rr_data_420,
        output wire [QNT_BIT-1:0] rr_data_421,
        output wire [QNT_BIT-1:0] rr_data_422,
        output wire [QNT_BIT-1:0] rr_data_423,
        output wire [QNT_BIT-1:0] rr_data_424,
        output wire [QNT_BIT-1:0] rr_data_425,
        output wire [QNT_BIT-1:0] rr_data_426,
        output wire [QNT_BIT-1:0] rr_data_427,
        output wire [QNT_BIT-1:0] rr_data_428,
        output wire [QNT_BIT-1:0] rr_data_429,
        output wire [QNT_BIT-1:0] rr_data_430,
        output wire [QNT_BIT-1:0] rr_data_431,
        output wire [QNT_BIT-1:0] rr_data_432,
        output wire [QNT_BIT-1:0] rr_data_433,
        output wire [QNT_BIT-1:0] rr_data_434,
        output wire [QNT_BIT-1:0] rr_data_435,
        output wire [QNT_BIT-1:0] rr_data_436,
        output wire [QNT_BIT-1:0] rr_data_437,
        output wire [QNT_BIT-1:0] rr_data_438,
        output wire [QNT_BIT-1:0] rr_data_439,
        output wire [QNT_BIT-1:0] rr_data_440,
        output wire [QNT_BIT-1:0] rr_data_441,
        output wire [QNT_BIT-1:0] rr_data_442,
        output wire [QNT_BIT-1:0] rr_data_443,
        output wire [QNT_BIT-1:0] rr_data_444,
        output wire [QNT_BIT-1:0] rr_data_445,
        output wire [QNT_BIT-1:0] rr_data_446,
        output wire [QNT_BIT-1:0] rr_data_447,
        output wire [QNT_BIT-1:0] rr_data_448,
        output wire [QNT_BIT-1:0] rr_data_449,
        output wire [QNT_BIT-1:0] rr_data_450,
        output wire [QNT_BIT-1:0] rr_data_451,
        output wire [QNT_BIT-1:0] rr_data_452,
        output wire [QNT_BIT-1:0] rr_data_453,
        output wire [QNT_BIT-1:0] rr_data_454,
        output wire [QNT_BIT-1:0] rr_data_455,
        output wire [QNT_BIT-1:0] rr_data_456,
        output wire [QNT_BIT-1:0] rr_data_457,
        output wire [QNT_BIT-1:0] rr_data_458,
        output wire [QNT_BIT-1:0] rr_data_459,
        output wire [QNT_BIT-1:0] rr_data_460,
        output wire [QNT_BIT-1:0] rr_data_461,
        output wire [QNT_BIT-1:0] rr_data_462,
        output wire [QNT_BIT-1:0] rr_data_463,
        output wire [QNT_BIT-1:0] rr_data_464,
        output wire [QNT_BIT-1:0] rr_data_465,
        output wire [QNT_BIT-1:0] rr_data_466,
        output wire [QNT_BIT-1:0] rr_data_467,
        output wire [QNT_BIT-1:0] rr_data_468,
        output wire [QNT_BIT-1:0] rr_data_469,
        output wire [QNT_BIT-1:0] rr_data_470,
        output wire [QNT_BIT-1:0] rr_data_471,
        output wire [QNT_BIT-1:0] rr_data_472,
        output wire [QNT_BIT-1:0] rr_data_473,
        output wire [QNT_BIT-1:0] rr_data_474,
        output wire [QNT_BIT-1:0] rr_data_475,
        output wire [QNT_BIT-1:0] rr_data_476,
        output wire [QNT_BIT-1:0] rr_data_477,
        output wire [QNT_BIT-1:0] rr_data_478,
        output wire [QNT_BIT-1:0] rr_data_479,
        output wire [QNT_BIT-1:0] rr_data_480,
        output wire [QNT_BIT-1:0] rr_data_481,
        output wire [QNT_BIT-1:0] rr_data_482,
        output wire [QNT_BIT-1:0] rr_data_483,
        output wire [QNT_BIT-1:0] rr_data_484,
        output wire [QNT_BIT-1:0] rr_data_485,
        output wire [QNT_BIT-1:0] rr_data_486,
        output wire [QNT_BIT-1:0] rr_data_487,
        output wire [QNT_BIT-1:0] rr_data_488,
        output wire [QNT_BIT-1:0] rr_data_489,
        output wire [QNT_BIT-1:0] rr_data_490,
        output wire [QNT_BIT-1:0] rr_data_491,
        output wire [QNT_BIT-1:0] rr_data_492,
        output wire [QNT_BIT-1:0] rr_data_493,
        output wire [QNT_BIT-1:0] rr_data_494,
        output wire [QNT_BIT-1:0] rr_data_495,
        output wire [QNT_BIT-1:0] rr_data_496,
        output wire [QNT_BIT-1:0] rr_data_497,
        output wire [QNT_BIT-1:0] rr_data_498,
        output wire [QNT_BIT-1:0] rr_data_499,
        output wire [QNT_BIT-1:0] rr_data_500,
        output wire [QNT_BIT-1:0] rr_data_501,
        output wire [QNT_BIT-1:0] rr_data_502,
        output wire [QNT_BIT-1:0] rr_data_503,
        output wire [QNT_BIT-1:0] rr_data_504,
        output wire [QNT_BIT-1:0] rr_data_505,
        output wire [QNT_BIT-1:0] rr_data_506,
        output wire [QNT_BIT-1:0] rr_data_507,
        output wire [QNT_BIT-1:0] rr_data_508,
        output wire [QNT_BIT-1:0] rr_data_509,
        output wire [QNT_BIT-1:0] rr_data_510,
        output wire [QNT_BIT-1:0] rr_data_511,
        output wire [QNT_BIT-1:0] rr_data_512,
        output wire [QNT_BIT-1:0] rr_data_513,
        output wire [QNT_BIT-1:0] rr_data_514,
        output wire [QNT_BIT-1:0] rr_data_515,
        output wire [QNT_BIT-1:0] rr_data_516,
        output wire [QNT_BIT-1:0] rr_data_517,
        output wire [QNT_BIT-1:0] rr_data_518,
        output wire [QNT_BIT-1:0] rr_data_519,
        output wire [QNT_BIT-1:0] rr_data_520,
        output wire [QNT_BIT-1:0] rr_data_521,
        output wire [QNT_BIT-1:0] rr_data_522,
        output wire [QNT_BIT-1:0] rr_data_523,
        output wire [QNT_BIT-1:0] rr_data_524,
        output wire [QNT_BIT-1:0] rr_data_525,
        output wire [QNT_BIT-1:0] rr_data_526,
        output wire [QNT_BIT-1:0] rr_data_527,
        output wire [QNT_BIT-1:0] rr_data_528,
        output wire [QNT_BIT-1:0] rr_data_529,
        output wire [QNT_BIT-1:0] rr_data_530,
        output wire [QNT_BIT-1:0] rr_data_531,
        output wire [QNT_BIT-1:0] rr_data_532,
        output wire [QNT_BIT-1:0] rr_data_533,
        output reg  [        6:0] addr,            // 写入 ram_llr 的内部地址
        output reg  [        1:0] flag_buffer_in,  // buffer 存有几帧信号
        output wire               flag_org_write_end,
        output wire               buffer_full      // 满了
    );

    // * 本文件主要是用来实现 buffer 的，重点在于生成地址信息和打一拍的写入数据
    // * 写入：采用乒乓操作。可以连续的读写
    // * 读出：对所有 24 个 combine_ram_llr 单元并行写入，所以只需要 24 个周期即可

    reg               write_en;  // 为 1 表示在输入数据过程中
    reg               write_en_reg;  // 多打一拍
    wire              write_page;  // 写入的 page 地址
    reg [9:0] write_col_cnt;  // 写入的 col 地址
    reg [6:0] write_cnt;  // 写入的单位矩阵内的地址
    reg [QNT_BIT-1:0] sink_reg;  // 打一拍和控制信号同步

    wire              read_page;  // 读取的 page 地址
    reg               read_en;
    reg [6:0] read_cnt;
    reg               read_end; // buffer 数据读取完成

    //************************************************************
    //*                       状态定义                           *
    //************************************************************
    localparam [2:0] IDLE = 3'b00_0;
    localparam [2:0] P0_write_P1_idle = 3'b10_0;
    localparam [2:0] P0_read_P1_write = 3'b11_1;
    localparam [2:0] P0_idle_P1_write = 3'b01_0;
    localparam [2:0] P0_write_P1_read = 3'b11_0;

    reg [2:0] current_state;
    reg [2:0] next_state;

    //************************************************************
    //*                       写逻辑                             *
    //************************************************************
    // 写入 en
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            write_en <= 1'b0;
        else if (sink_star == 1'b1 && !buffer_full)
            write_en <= 1'b1;
        else if (sink_stop == 1'b1)
            write_en <= 1'b0;
        else
            write_en <= write_en;


    // 多打一拍 reg
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            write_en_reg <= 1'b0;
        else
            write_en_reg <= write_en;


    // 生成写入的单位矩阵内的地址
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            write_cnt <= 7'b0;
        else if (write_cnt == QC_LDPC_BLOCK_SIZE - 1 || sink_stop == 1'b1)
            write_cnt <= 7'b0;
        else if (write_en == 1'b1)
            write_cnt <= write_cnt + 1'b1;
        else
            write_cnt <= write_cnt;


    // 生成写入的 col 地址
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            write_col_cnt <= 10'b0;
        else if ((write_col_cnt == QC_LDPC_COL_COUNT - 1 && write_cnt == QC_LDPC_BLOCK_SIZE - 1) || sink_star == 1'b1)
            write_col_cnt <= 10'b0;
        else if (write_cnt == QC_LDPC_BLOCK_SIZE - 1)
            write_col_cnt <= write_col_cnt + 1'b1;
        else
            write_col_cnt <= write_col_cnt;


    // 写入页地址，用 wire 以实现时序对齐
    assign write_page = (current_state == P0_read_P1_write) || (current_state == P0_idle_P1_write);


    // 存有帧的个数
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            flag_buffer_in <= 2'b0;
        else if ((write_en_reg == 1'b1 && sink_stop == 1'b1) && read_end == 1'b1)
            flag_buffer_in <= flag_buffer_in;
        else if (write_en_reg == 1'b1 && sink_stop == 1'b1) // 存入一帧
            flag_buffer_in <= flag_buffer_in + 2'b1;
        else if (read_end == 1'b1) // 读完一帧
            flag_buffer_in <= flag_buffer_in - 2'b1;
        else 
            flag_buffer_in <= flag_buffer_in;


    // 写满信号
    assign buffer_full = (current_state == P0_read_P1_write) || (current_state == P0_write_P1_read);


    // 打一拍 sink
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            sink_reg <= 1'b0;
        else
            sink_reg <= sink;


    //************************************************************
    //*                       读逻辑                              *
    //************************************************************
    // 读 en
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            read_en <= 1'b0;
        else if (flag_org_update == 1'b1)
            read_en <= 1'b1;
        else if (read_cnt == QC_LDPC_BLOCK_SIZE - 1)
            read_en <= 1'b0;
        else
            read_en <= read_en;


    // 读 end
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            read_end <= 1'b0;
        else if (read_cnt == QC_LDPC_BLOCK_SIZE - 1)
            read_end <= 1'b1;
        else
            read_end <= 1'b0;


    // 生成写入的单位矩阵内的地址
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            read_cnt <= 8'b0;
        else if (read_cnt == QC_LDPC_BLOCK_SIZE - 1)
            read_cnt <= 8'b0;
        else if (read_en == 1'b1)
            read_cnt <= read_cnt + 1'b1;
        else
            read_cnt <= read_cnt;


    // 读页地址
    assign read_page = (current_state == P0_idle_P1_write) || (current_state == P0_write_P1_read);


    // 打一拍的 en 输出，等待 ram 读的一个周期延迟
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n  == 1'b0)
            buffer_wr_en <= 1'b0;
        else
            buffer_wr_en <= read_en;


    // 打一拍的 addr 输出，等待 ram 读的一个周期延迟
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n  == 1'b0)
            addr <= 8'b0;
        else
            addr <= read_cnt;


    assign flag_org_write_end = read_end;

    //************************************************************
    //*                       状态机                             *
    //************************************************************
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            current_state <= IDLE;  // 复位时回到IDLE状态
        else
            current_state <= next_state;  // 否则更新到下一状态


    always @(*)
    case (current_state)
        IDLE: begin
            if (sink_star)
                next_state = P0_write_P1_idle;
            else
                next_state = next_state;
        end
        P0_write_P1_idle: begin
            if (sink_star && read_end)
                next_state = next_state;
            else if (sink_star)
                next_state = P0_read_P1_write;
            else if (read_end)
                next_state = IDLE;
            else
                next_state = next_state;
        end
        P0_read_P1_write: begin
            if (read_end)
                next_state = P0_idle_P1_write;
            else
                next_state = next_state;
        end
        P0_idle_P1_write: begin
            if (sink_star && read_end)
                next_state = next_state;
            else if (sink_star)
                next_state = P0_write_P1_read;
            else if (read_end)
                next_state = IDLE;
            else
                next_state = next_state;
        end
        P0_write_P1_read: begin
            if (read_end)
                next_state = P0_write_P1_idle;
            else
                next_state = next_state;
        end
        default:
            next_state = IDLE;
    endcase


    //************************************************************
    //*                       实例化                              *
    //************************************************************

    buffer_ram #(
                   .QNT_BIT           (QNT_BIT),
                   .QC_LDPC_COL_COUNT (QC_LDPC_COL_COUNT),
                   .QC_LDPC_BLOCK_SIZE(QC_LDPC_BLOCK_SIZE)
               ) u_buffer_ram (
                   .sys_clk      (sys_clk),
                   .sys_rst_n    (sys_rst_n),
                   .write_en     (write_en),
                   .write_page   (write_page),
                   .write_col_cnt(write_col_cnt),
                   .write_cnt    (write_cnt),
                   .sink         (sink_reg),
                   .read_en      (read_en),
                   .read_page    (read_page),
                   .read_cnt     (read_cnt),

                   .rr_data_1 (rr_data_1),
                   .rr_data_2 (rr_data_2),
                   .rr_data_3 (rr_data_3),
                   .rr_data_4 (rr_data_4),
                   .rr_data_5 (rr_data_5),
                   .rr_data_6 (rr_data_6),
                   .rr_data_7 (rr_data_7),
                   .rr_data_8 (rr_data_8),
                   .rr_data_9 (rr_data_9),
                   .rr_data_10(rr_data_10),
                   .rr_data_11(rr_data_11),
                   .rr_data_12(rr_data_12),
                   .rr_data_13(rr_data_13),
                   .rr_data_14(rr_data_14),
                   .rr_data_15(rr_data_15),
                   .rr_data_16(rr_data_16),
                   .rr_data_17(rr_data_17),
                   .rr_data_18(rr_data_18),
                   .rr_data_19(rr_data_19),
                   .rr_data_20(rr_data_20),
                   .rr_data_21(rr_data_21),
                   .rr_data_22(rr_data_22),
                   .rr_data_23(rr_data_23),
                   .rr_data_24(rr_data_24),
                   .rr_data_25(rr_data_25),
                   .rr_data_26(rr_data_26),
                   .rr_data_27(rr_data_27),
                   .rr_data_28(rr_data_28),
                   .rr_data_29(rr_data_29),
                   .rr_data_30(rr_data_30),
                   .rr_data_31(rr_data_31),
                   .rr_data_32(rr_data_32),
                   .rr_data_33(rr_data_33),
                   .rr_data_34(rr_data_34),
                   .rr_data_35(rr_data_35),
                   .rr_data_36(rr_data_36),
                   .rr_data_37(rr_data_37),
                   .rr_data_38(rr_data_38),
                   .rr_data_39(rr_data_39),
                   .rr_data_40(rr_data_40),
                   .rr_data_41(rr_data_41),
                   .rr_data_42(rr_data_42),
                   .rr_data_43(rr_data_43),
                   .rr_data_44(rr_data_44),
                   .rr_data_45(rr_data_45),
                   .rr_data_46(rr_data_46),
                   .rr_data_47(rr_data_47),
                   .rr_data_48(rr_data_48),
                   .rr_data_49(rr_data_49),
                   .rr_data_50(rr_data_50),
                   .rr_data_51(rr_data_51),
                   .rr_data_52(rr_data_52),
                   .rr_data_53(rr_data_53),
                   .rr_data_54(rr_data_54),
                   .rr_data_55(rr_data_55),
                   .rr_data_56(rr_data_56),
                   .rr_data_57(rr_data_57),
                   .rr_data_58(rr_data_58),
                   .rr_data_59(rr_data_59),
                   .rr_data_60(rr_data_60),
                   .rr_data_61(rr_data_61),
                   .rr_data_62(rr_data_62),
                   .rr_data_63(rr_data_63),
                   .rr_data_64(rr_data_64),
                   .rr_data_65(rr_data_65),
                   .rr_data_66(rr_data_66),
                   .rr_data_67(rr_data_67),
                   .rr_data_68(rr_data_68),
                   .rr_data_69(rr_data_69),
                   .rr_data_70(rr_data_70),
                   .rr_data_71(rr_data_71),
                   .rr_data_72(rr_data_72),
                   .rr_data_73(rr_data_73),
                   .rr_data_74(rr_data_74),
                   .rr_data_75(rr_data_75),
                   .rr_data_76(rr_data_76),
                   .rr_data_77(rr_data_77),
                   .rr_data_78(rr_data_78),
                   .rr_data_79(rr_data_79),
                   .rr_data_80(rr_data_80),
                   .rr_data_81(rr_data_81),
                   .rr_data_82(rr_data_82),
                   .rr_data_83(rr_data_83),
                   .rr_data_84(rr_data_84),
                   .rr_data_85(rr_data_85),
                   .rr_data_86(rr_data_86),
                   .rr_data_87(rr_data_87),
                   .rr_data_88(rr_data_88),
                   .rr_data_89(rr_data_89),
                   .rr_data_90(rr_data_90),
                   .rr_data_91(rr_data_91),
                   .rr_data_92(rr_data_92),
                   .rr_data_93(rr_data_93),
                   .rr_data_94(rr_data_94),
                   .rr_data_95(rr_data_95),
                   .rr_data_96(rr_data_96),
                   .rr_data_97(rr_data_97),
                   .rr_data_98(rr_data_98),
                   .rr_data_99(rr_data_99),
                   .rr_data_100(rr_data_100),
                   .rr_data_101(rr_data_101),
                   .rr_data_102(rr_data_102),
                   .rr_data_103(rr_data_103),
                   .rr_data_104(rr_data_104),
                   .rr_data_105(rr_data_105),
                   .rr_data_106(rr_data_106),
                   .rr_data_107(rr_data_107),
                   .rr_data_108(rr_data_108),
                   .rr_data_109(rr_data_109),
                   .rr_data_110(rr_data_110),
                   .rr_data_111(rr_data_111),
                   .rr_data_112(rr_data_112),
                   .rr_data_113(rr_data_113),
                   .rr_data_114(rr_data_114),
                   .rr_data_115(rr_data_115),
                   .rr_data_116(rr_data_116),
                   .rr_data_117(rr_data_117),
                   .rr_data_118(rr_data_118),
                   .rr_data_119(rr_data_119),
                   .rr_data_120(rr_data_120),
                   .rr_data_121(rr_data_121),
                   .rr_data_122(rr_data_122),
                   .rr_data_123(rr_data_123),
                   .rr_data_124(rr_data_124),
                   .rr_data_125(rr_data_125),
                   .rr_data_126(rr_data_126),
                   .rr_data_127(rr_data_127),
                   .rr_data_128(rr_data_128),
                   .rr_data_129(rr_data_129),
                   .rr_data_130(rr_data_130),
                   .rr_data_131(rr_data_131),
                   .rr_data_132(rr_data_132),
                   .rr_data_133(rr_data_133),
                   .rr_data_134(rr_data_134),
                   .rr_data_135(rr_data_135),
                   .rr_data_136(rr_data_136),
                   .rr_data_137(rr_data_137),
                   .rr_data_138(rr_data_138),
                   .rr_data_139(rr_data_139),
                   .rr_data_140(rr_data_140),
                   .rr_data_141(rr_data_141),
                   .rr_data_142(rr_data_142),
                   .rr_data_143(rr_data_143),
                   .rr_data_144(rr_data_144),
                   .rr_data_145(rr_data_145),
                   .rr_data_146(rr_data_146),
                   .rr_data_147(rr_data_147),
                   .rr_data_148(rr_data_148),
                   .rr_data_149(rr_data_149),
                   .rr_data_150(rr_data_150),
                   .rr_data_151(rr_data_151),
                   .rr_data_152(rr_data_152),
                   .rr_data_153(rr_data_153),
                   .rr_data_154(rr_data_154),
                   .rr_data_155(rr_data_155),
                   .rr_data_156(rr_data_156),
                   .rr_data_157(rr_data_157),
                   .rr_data_158(rr_data_158),
                   .rr_data_159(rr_data_159),
                   .rr_data_160(rr_data_160),
                   .rr_data_161(rr_data_161),
                   .rr_data_162(rr_data_162),
                   .rr_data_163(rr_data_163),
                   .rr_data_164(rr_data_164),
                   .rr_data_165(rr_data_165),
                   .rr_data_166(rr_data_166),
                   .rr_data_167(rr_data_167),
                   .rr_data_168(rr_data_168),
                   .rr_data_169(rr_data_169),
                   .rr_data_170(rr_data_170),
                   .rr_data_171(rr_data_171),
                   .rr_data_172(rr_data_172),
                   .rr_data_173(rr_data_173),
                   .rr_data_174(rr_data_174),
                   .rr_data_175(rr_data_175),
                   .rr_data_176(rr_data_176),
                   .rr_data_177(rr_data_177),
                   .rr_data_178(rr_data_178),
                   .rr_data_179(rr_data_179),
                   .rr_data_180(rr_data_180),
                   .rr_data_181(rr_data_181),
                   .rr_data_182(rr_data_182),
                   .rr_data_183(rr_data_183),
                   .rr_data_184(rr_data_184),
                   .rr_data_185(rr_data_185),
                   .rr_data_186(rr_data_186),
                   .rr_data_187(rr_data_187),
                   .rr_data_188(rr_data_188),
                   .rr_data_189(rr_data_189),
                   .rr_data_190(rr_data_190),
                   .rr_data_191(rr_data_191),
                   .rr_data_192(rr_data_192),
                   .rr_data_193(rr_data_193),
                   .rr_data_194(rr_data_194),
                   .rr_data_195(rr_data_195),
                   .rr_data_196(rr_data_196),
                   .rr_data_197(rr_data_197),
                   .rr_data_198(rr_data_198),
                   .rr_data_199(rr_data_199),
                   .rr_data_200(rr_data_200),
                   .rr_data_201(rr_data_201),
                   .rr_data_202(rr_data_202),
                   .rr_data_203(rr_data_203),
                   .rr_data_204(rr_data_204),
                   .rr_data_205(rr_data_205),
                   .rr_data_206(rr_data_206),
                   .rr_data_207(rr_data_207),
                   .rr_data_208(rr_data_208),
                   .rr_data_209(rr_data_209),
                   .rr_data_210(rr_data_210),
                   .rr_data_211(rr_data_211),
                   .rr_data_212(rr_data_212),
                   .rr_data_213(rr_data_213),
                   .rr_data_214(rr_data_214),
                   .rr_data_215(rr_data_215),
                   .rr_data_216(rr_data_216),
                   .rr_data_217(rr_data_217),
                   .rr_data_218(rr_data_218),
                   .rr_data_219(rr_data_219),
                   .rr_data_220(rr_data_220),
                   .rr_data_221(rr_data_221),
                   .rr_data_222(rr_data_222),
                   .rr_data_223(rr_data_223),
                   .rr_data_224(rr_data_224),
                   .rr_data_225(rr_data_225),
                   .rr_data_226(rr_data_226),
                   .rr_data_227(rr_data_227),
                   .rr_data_228(rr_data_228),
                   .rr_data_229(rr_data_229),
                   .rr_data_230(rr_data_230),
                   .rr_data_231(rr_data_231),
                   .rr_data_232(rr_data_232),
                   .rr_data_233(rr_data_233),
                   .rr_data_234(rr_data_234),
                   .rr_data_235(rr_data_235),
                   .rr_data_236(rr_data_236),
                   .rr_data_237(rr_data_237),
                   .rr_data_238(rr_data_238),
                   .rr_data_239(rr_data_239),
                   .rr_data_240(rr_data_240),
                   .rr_data_241(rr_data_241),
                   .rr_data_242(rr_data_242),
                   .rr_data_243(rr_data_243),
                   .rr_data_244(rr_data_244),
                   .rr_data_245(rr_data_245),
                   .rr_data_246(rr_data_246),
                   .rr_data_247(rr_data_247),
                   .rr_data_248(rr_data_248),
                   .rr_data_249(rr_data_249),
                   .rr_data_250(rr_data_250),
                   .rr_data_251(rr_data_251),
                   .rr_data_252(rr_data_252),
                   .rr_data_253(rr_data_253),
                   .rr_data_254(rr_data_254),
                   .rr_data_255(rr_data_255),
                   .rr_data_256(rr_data_256),
                   .rr_data_257(rr_data_257),
                   .rr_data_258(rr_data_258),
                   .rr_data_259(rr_data_259),
                   .rr_data_260(rr_data_260),
                   .rr_data_261(rr_data_261),
                   .rr_data_262(rr_data_262),
                   .rr_data_263(rr_data_263),
                   .rr_data_264(rr_data_264),
                   .rr_data_265(rr_data_265),
                   .rr_data_266(rr_data_266),
                   .rr_data_267(rr_data_267),
                   .rr_data_268(rr_data_268),
                   .rr_data_269(rr_data_269),
                   .rr_data_270(rr_data_270),
                   .rr_data_271(rr_data_271),
                   .rr_data_272(rr_data_272),
                   .rr_data_273(rr_data_273),
                   .rr_data_274(rr_data_274),
                   .rr_data_275(rr_data_275),
                   .rr_data_276(rr_data_276),
                   .rr_data_277(rr_data_277),
                   .rr_data_278(rr_data_278),
                   .rr_data_279(rr_data_279),
                   .rr_data_280(rr_data_280),
                   .rr_data_281(rr_data_281),
                   .rr_data_282(rr_data_282),
                   .rr_data_283(rr_data_283),
                   .rr_data_284(rr_data_284),
                   .rr_data_285(rr_data_285),
                   .rr_data_286(rr_data_286),
                   .rr_data_287(rr_data_287),
                   .rr_data_288(rr_data_288),
                   .rr_data_289(rr_data_289),
                   .rr_data_290(rr_data_290),
                   .rr_data_291(rr_data_291),
                   .rr_data_292(rr_data_292),
                   .rr_data_293(rr_data_293),
                   .rr_data_294(rr_data_294),
                   .rr_data_295(rr_data_295),
                   .rr_data_296(rr_data_296),
                   .rr_data_297(rr_data_297),
                   .rr_data_298(rr_data_298),
                   .rr_data_299(rr_data_299),
                   .rr_data_300(rr_data_300),
                   .rr_data_301(rr_data_301),
                   .rr_data_302(rr_data_302),
                   .rr_data_303(rr_data_303),
                   .rr_data_304(rr_data_304),
                   .rr_data_305(rr_data_305),
                   .rr_data_306(rr_data_306),
                   .rr_data_307(rr_data_307),
                   .rr_data_308(rr_data_308),
                   .rr_data_309(rr_data_309),
                   .rr_data_310(rr_data_310),
                   .rr_data_311(rr_data_311),
                   .rr_data_312(rr_data_312),
                   .rr_data_313(rr_data_313),
                   .rr_data_314(rr_data_314),
                   .rr_data_315(rr_data_315),
                   .rr_data_316(rr_data_316),
                   .rr_data_317(rr_data_317),
                   .rr_data_318(rr_data_318),
                   .rr_data_319(rr_data_319),
                   .rr_data_320(rr_data_320),
                   .rr_data_321(rr_data_321),
                   .rr_data_322(rr_data_322),
                   .rr_data_323(rr_data_323),
                   .rr_data_324(rr_data_324),
                   .rr_data_325(rr_data_325),
                   .rr_data_326(rr_data_326),
                   .rr_data_327(rr_data_327),
                   .rr_data_328(rr_data_328),
                   .rr_data_329(rr_data_329),
                   .rr_data_330(rr_data_330),
                   .rr_data_331(rr_data_331),
                   .rr_data_332(rr_data_332),
                   .rr_data_333(rr_data_333),
                   .rr_data_334(rr_data_334),
                   .rr_data_335(rr_data_335),
                   .rr_data_336(rr_data_336),
                   .rr_data_337(rr_data_337),
                   .rr_data_338(rr_data_338),
                   .rr_data_339(rr_data_339),
                   .rr_data_340(rr_data_340),
                   .rr_data_341(rr_data_341),
                   .rr_data_342(rr_data_342),
                   .rr_data_343(rr_data_343),
                   .rr_data_344(rr_data_344),
                   .rr_data_345(rr_data_345),
                   .rr_data_346(rr_data_346),
                   .rr_data_347(rr_data_347),
                   .rr_data_348(rr_data_348),
                   .rr_data_349(rr_data_349),
                   .rr_data_350(rr_data_350),
                   .rr_data_351(rr_data_351),
                   .rr_data_352(rr_data_352),
                   .rr_data_353(rr_data_353),
                   .rr_data_354(rr_data_354),
                   .rr_data_355(rr_data_355),
                   .rr_data_356(rr_data_356),
                   .rr_data_357(rr_data_357),
                   .rr_data_358(rr_data_358),
                   .rr_data_359(rr_data_359),
                   .rr_data_360(rr_data_360),
                   .rr_data_361(rr_data_361),
                   .rr_data_362(rr_data_362),
                   .rr_data_363(rr_data_363),
                   .rr_data_364(rr_data_364),
                   .rr_data_365(rr_data_365),
                   .rr_data_366(rr_data_366),
                   .rr_data_367(rr_data_367),
                   .rr_data_368(rr_data_368),
                   .rr_data_369(rr_data_369),
                   .rr_data_370(rr_data_370),
                   .rr_data_371(rr_data_371),
                   .rr_data_372(rr_data_372),
                   .rr_data_373(rr_data_373),
                   .rr_data_374(rr_data_374),
                   .rr_data_375(rr_data_375),
                   .rr_data_376(rr_data_376),
                   .rr_data_377(rr_data_377),
                   .rr_data_378(rr_data_378),
                   .rr_data_379(rr_data_379),
                   .rr_data_380(rr_data_380),
                   .rr_data_381(rr_data_381),
                   .rr_data_382(rr_data_382),
                   .rr_data_383(rr_data_383),
                   .rr_data_384(rr_data_384),
                   .rr_data_385(rr_data_385),
                   .rr_data_386(rr_data_386),
                   .rr_data_387(rr_data_387),
                   .rr_data_388(rr_data_388),
                   .rr_data_389(rr_data_389),
                   .rr_data_390(rr_data_390),
                   .rr_data_391(rr_data_391),
                   .rr_data_392(rr_data_392),
                   .rr_data_393(rr_data_393),
                   .rr_data_394(rr_data_394),
                   .rr_data_395(rr_data_395),
                   .rr_data_396(rr_data_396),
                   .rr_data_397(rr_data_397),
                   .rr_data_398(rr_data_398),
                   .rr_data_399(rr_data_399),
                   .rr_data_400(rr_data_400),
                   .rr_data_401(rr_data_401),
                   .rr_data_402(rr_data_402),
                   .rr_data_403(rr_data_403),
                   .rr_data_404(rr_data_404),
                   .rr_data_405(rr_data_405),
                   .rr_data_406(rr_data_406),
                   .rr_data_407(rr_data_407),
                   .rr_data_408(rr_data_408),
                   .rr_data_409(rr_data_409),
                   .rr_data_410(rr_data_410),
                   .rr_data_411(rr_data_411),
                   .rr_data_412(rr_data_412),
                   .rr_data_413(rr_data_413),
                   .rr_data_414(rr_data_414),
                   .rr_data_415(rr_data_415),
                   .rr_data_416(rr_data_416),
                   .rr_data_417(rr_data_417),
                   .rr_data_418(rr_data_418),
                   .rr_data_419(rr_data_419),
                   .rr_data_420(rr_data_420),
                   .rr_data_421(rr_data_421),
                   .rr_data_422(rr_data_422),
                   .rr_data_423(rr_data_423),
                   .rr_data_424(rr_data_424),
                   .rr_data_425(rr_data_425),
                   .rr_data_426(rr_data_426),
                   .rr_data_427(rr_data_427),
                   .rr_data_428(rr_data_428),
                   .rr_data_429(rr_data_429),
                   .rr_data_430(rr_data_430),
                   .rr_data_431(rr_data_431),
                   .rr_data_432(rr_data_432),
                   .rr_data_433(rr_data_433),
                   .rr_data_434(rr_data_434),
                   .rr_data_435(rr_data_435),
                   .rr_data_436(rr_data_436),
                   .rr_data_437(rr_data_437),
                   .rr_data_438(rr_data_438),
                   .rr_data_439(rr_data_439),
                   .rr_data_440(rr_data_440),
                   .rr_data_441(rr_data_441),
                   .rr_data_442(rr_data_442),
                   .rr_data_443(rr_data_443),
                   .rr_data_444(rr_data_444),
                   .rr_data_445(rr_data_445),
                   .rr_data_446(rr_data_446),
                   .rr_data_447(rr_data_447),
                   .rr_data_448(rr_data_448),
                   .rr_data_449(rr_data_449),
                   .rr_data_450(rr_data_450),
                   .rr_data_451(rr_data_451),
                   .rr_data_452(rr_data_452),
                   .rr_data_453(rr_data_453),
                   .rr_data_454(rr_data_454),
                   .rr_data_455(rr_data_455),
                   .rr_data_456(rr_data_456),
                   .rr_data_457(rr_data_457),
                   .rr_data_458(rr_data_458),
                   .rr_data_459(rr_data_459),
                   .rr_data_460(rr_data_460),
                   .rr_data_461(rr_data_461),
                   .rr_data_462(rr_data_462),
                   .rr_data_463(rr_data_463),
                   .rr_data_464(rr_data_464),
                   .rr_data_465(rr_data_465),
                   .rr_data_466(rr_data_466),
                   .rr_data_467(rr_data_467),
                   .rr_data_468(rr_data_468),
                   .rr_data_469(rr_data_469),
                   .rr_data_470(rr_data_470),
                   .rr_data_471(rr_data_471),
                   .rr_data_472(rr_data_472),
                   .rr_data_473(rr_data_473),
                   .rr_data_474(rr_data_474),
                   .rr_data_475(rr_data_475),
                   .rr_data_476(rr_data_476),
                   .rr_data_477(rr_data_477),
                   .rr_data_478(rr_data_478),
                   .rr_data_479(rr_data_479),
                   .rr_data_480(rr_data_480),
                   .rr_data_481(rr_data_481),
                   .rr_data_482(rr_data_482),
                   .rr_data_483(rr_data_483),
                   .rr_data_484(rr_data_484),
                   .rr_data_485(rr_data_485),
                   .rr_data_486(rr_data_486),
                   .rr_data_487(rr_data_487),
                   .rr_data_488(rr_data_488),
                   .rr_data_489(rr_data_489),
                   .rr_data_490(rr_data_490),
                   .rr_data_491(rr_data_491),
                   .rr_data_492(rr_data_492),
                   .rr_data_493(rr_data_493),
                   .rr_data_494(rr_data_494),
                   .rr_data_495(rr_data_495),
                   .rr_data_496(rr_data_496),
                   .rr_data_497(rr_data_497),
                   .rr_data_498(rr_data_498),
                   .rr_data_499(rr_data_499),
                   .rr_data_500(rr_data_500),
                   .rr_data_501(rr_data_501),
                   .rr_data_502(rr_data_502),
                   .rr_data_503(rr_data_503),
                   .rr_data_504(rr_data_504),
                   .rr_data_505(rr_data_505),
                   .rr_data_506(rr_data_506),
                   .rr_data_507(rr_data_507),
                   .rr_data_508(rr_data_508),
                   .rr_data_509(rr_data_509),
                   .rr_data_510(rr_data_510),
                   .rr_data_511(rr_data_511),
                   .rr_data_512(rr_data_512),
                   .rr_data_513(rr_data_513),
                   .rr_data_514(rr_data_514),
                   .rr_data_515(rr_data_515),
                   .rr_data_516(rr_data_516),
                   .rr_data_517(rr_data_517),
                   .rr_data_518(rr_data_518),
                   .rr_data_519(rr_data_519),
                   .rr_data_520(rr_data_520),
                   .rr_data_521(rr_data_521),
                   .rr_data_522(rr_data_522),
                   .rr_data_523(rr_data_523),
                   .rr_data_524(rr_data_524),
                   .rr_data_525(rr_data_525),
                   .rr_data_526(rr_data_526),
                   .rr_data_527(rr_data_527),
                   .rr_data_528(rr_data_528),
                   .rr_data_529(rr_data_529),
                   .rr_data_530(rr_data_530),
                   .rr_data_531(rr_data_531),
                   .rr_data_532(rr_data_532),
                   .rr_data_533(rr_data_533)
               );

endmodule
