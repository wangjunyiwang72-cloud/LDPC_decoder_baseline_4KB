module buffer_ram #(
        parameter QNT_BIT            = 4,  // LLR量化位宽4位
        parameter QC_LDPC_COL_COUNT  = 533,  // 基矩阵列数
        parameter QC_LDPC_BLOCK_SIZE = 64   // 扩展因子
    ) (
        input wire sys_clk,
        input wire sys_rst_n,

        // 写通道
        input wire               write_en,       // 写有效信号
        input wire               write_page,     // 写入的 page 地址
        input wire [9:0] write_col_cnt,  // 写入的 col 地址
        input wire [7:0] write_cnt,      // 写入的单位矩阵内的地址
        input wire [QNT_BIT-1:0] sink,           // 输入数据

        // 读通道
        input  wire               read_en,     // 读有效信号
        input  wire               read_page,   // 读取的 page 地址
        input  wire [7:0] read_cnt,    // 读取的单位矩阵内的地址
        output wire [QNT_BIT-1:0] rr_data_1,
        output wire [QNT_BIT-1:0] rr_data_2,
        output wire [QNT_BIT-1:0] rr_data_3,
        output wire [QNT_BIT-1:0] rr_data_4,
        output wire [QNT_BIT-1:0] rr_data_5,
        output wire [QNT_BIT-1:0] rr_data_6,
        output wire [QNT_BIT-1:0] rr_data_7,
        output wire [QNT_BIT-1:0] rr_data_8,
        output wire [QNT_BIT-1:0] rr_data_9,
        output wire [QNT_BIT-1:0] rr_data_10,
        output wire [QNT_BIT-1:0] rr_data_11,
        output wire [QNT_BIT-1:0] rr_data_12,
        output wire [QNT_BIT-1:0] rr_data_13,
        output wire [QNT_BIT-1:0] rr_data_14,
        output wire [QNT_BIT-1:0] rr_data_15,
        output wire [QNT_BIT-1:0] rr_data_16,
        output wire [QNT_BIT-1:0] rr_data_17,
        output wire [QNT_BIT-1:0] rr_data_18,
        output wire [QNT_BIT-1:0] rr_data_19,
        output wire [QNT_BIT-1:0] rr_data_20,
        output wire [QNT_BIT-1:0] rr_data_21,
        output wire [QNT_BIT-1:0] rr_data_22,
        output wire [QNT_BIT-1:0] rr_data_23,
        output wire [QNT_BIT-1:0] rr_data_24,
        output wire [QNT_BIT-1:0] rr_data_25,
        output wire [QNT_BIT-1:0] rr_data_26,
        output wire [QNT_BIT-1:0] rr_data_27,
        output wire [QNT_BIT-1:0] rr_data_28,
        output wire [QNT_BIT-1:0] rr_data_29,
        output wire [QNT_BIT-1:0] rr_data_30,
        output wire [QNT_BIT-1:0] rr_data_31,
        output wire [QNT_BIT-1:0] rr_data_32,
        output wire [QNT_BIT-1:0] rr_data_33,
        output wire [QNT_BIT-1:0] rr_data_34,
        output wire [QNT_BIT-1:0] rr_data_35,
        output wire [QNT_BIT-1:0] rr_data_36,
        output wire [QNT_BIT-1:0] rr_data_37,
        output wire [QNT_BIT-1:0] rr_data_38,
        output wire [QNT_BIT-1:0] rr_data_39,
        output wire [QNT_BIT-1:0] rr_data_40,
        output wire [QNT_BIT-1:0] rr_data_41,
        output wire [QNT_BIT-1:0] rr_data_42,
        output wire [QNT_BIT-1:0] rr_data_43,
        output wire [QNT_BIT-1:0] rr_data_44,
        output wire [QNT_BIT-1:0] rr_data_45,
        output wire [QNT_BIT-1:0] rr_data_46,
        output wire [QNT_BIT-1:0] rr_data_47,
        output wire [QNT_BIT-1:0] rr_data_48,
        output wire [QNT_BIT-1:0] rr_data_49,
        output wire [QNT_BIT-1:0] rr_data_50,
        output wire [QNT_BIT-1:0] rr_data_51,
        output wire [QNT_BIT-1:0] rr_data_52,
        output wire [QNT_BIT-1:0] rr_data_53,
        output wire [QNT_BIT-1:0] rr_data_54,
        output wire [QNT_BIT-1:0] rr_data_55,
        output wire [QNT_BIT-1:0] rr_data_56,
        output wire [QNT_BIT-1:0] rr_data_57,
        output wire [QNT_BIT-1:0] rr_data_58,
        output wire [QNT_BIT-1:0] rr_data_59,
        output wire [QNT_BIT-1:0] rr_data_60,
        output wire [QNT_BIT-1:0] rr_data_61,
        output wire [QNT_BIT-1:0] rr_data_62,
        output wire [QNT_BIT-1:0] rr_data_63,
        output wire [QNT_BIT-1:0] rr_data_64,
        output wire [QNT_BIT-1:0] rr_data_65,
        output wire [QNT_BIT-1:0] rr_data_66,
        output wire [QNT_BIT-1:0] rr_data_67,
        output wire [QNT_BIT-1:0] rr_data_68,
        output wire [QNT_BIT-1:0] rr_data_69,
        output wire [QNT_BIT-1:0] rr_data_70,
        output wire [QNT_BIT-1:0] rr_data_71,
        output wire [QNT_BIT-1:0] rr_data_72,
        output wire [QNT_BIT-1:0] rr_data_73,
        output wire [QNT_BIT-1:0] rr_data_74,
        output wire [QNT_BIT-1:0] rr_data_75,
        output wire [QNT_BIT-1:0] rr_data_76,
        output wire [QNT_BIT-1:0] rr_data_77,
        output wire [QNT_BIT-1:0] rr_data_78,
        output wire [QNT_BIT-1:0] rr_data_79,
        output wire [QNT_BIT-1:0] rr_data_80,
        output wire [QNT_BIT-1:0] rr_data_81,
        output wire [QNT_BIT-1:0] rr_data_82,
        output wire [QNT_BIT-1:0] rr_data_83,
        output wire [QNT_BIT-1:0] rr_data_84,
        output wire [QNT_BIT-1:0] rr_data_85,
        output wire [QNT_BIT-1:0] rr_data_86,
        output wire [QNT_BIT-1:0] rr_data_87,
        output wire [QNT_BIT-1:0] rr_data_88,
        output wire [QNT_BIT-1:0] rr_data_89,
        output wire [QNT_BIT-1:0] rr_data_90,
        output wire [QNT_BIT-1:0] rr_data_91,
        output wire [QNT_BIT-1:0] rr_data_92,
        output wire [QNT_BIT-1:0] rr_data_93,
        output wire [QNT_BIT-1:0] rr_data_94,
        output wire [QNT_BIT-1:0] rr_data_95,
        output wire [QNT_BIT-1:0] rr_data_96,
        output wire [QNT_BIT-1:0] rr_data_97,
        output wire [QNT_BIT-1:0] rr_data_98,
        output wire [QNT_BIT-1:0] rr_data_99,
        output wire [QNT_BIT-1:0] rr_data_100,
        output wire [QNT_BIT-1:0] rr_data_101,
        output wire [QNT_BIT-1:0] rr_data_102,
        output wire [QNT_BIT-1:0] rr_data_103,
        output wire [QNT_BIT-1:0] rr_data_104,
        output wire [QNT_BIT-1:0] rr_data_105,
        output wire [QNT_BIT-1:0] rr_data_106,
        output wire [QNT_BIT-1:0] rr_data_107,
        output wire [QNT_BIT-1:0] rr_data_108,
        output wire [QNT_BIT-1:0] rr_data_109,
        output wire [QNT_BIT-1:0] rr_data_110,
        output wire [QNT_BIT-1:0] rr_data_111,
        output wire [QNT_BIT-1:0] rr_data_112,
        output wire [QNT_BIT-1:0] rr_data_113,
        output wire [QNT_BIT-1:0] rr_data_114,
        output wire [QNT_BIT-1:0] rr_data_115,
        output wire [QNT_BIT-1:0] rr_data_116,
        output wire [QNT_BIT-1:0] rr_data_117,
        output wire [QNT_BIT-1:0] rr_data_118,
        output wire [QNT_BIT-1:0] rr_data_119,
        output wire [QNT_BIT-1:0] rr_data_120,
        output wire [QNT_BIT-1:0] rr_data_121,
        output wire [QNT_BIT-1:0] rr_data_122,
        output wire [QNT_BIT-1:0] rr_data_123,
        output wire [QNT_BIT-1:0] rr_data_124,
        output wire [QNT_BIT-1:0] rr_data_125,
        output wire [QNT_BIT-1:0] rr_data_126,
        output wire [QNT_BIT-1:0] rr_data_127,
        output wire [QNT_BIT-1:0] rr_data_128,
        output wire [QNT_BIT-1:0] rr_data_129,
        output wire [QNT_BIT-1:0] rr_data_130,
        output wire [QNT_BIT-1:0] rr_data_131,
        output wire [QNT_BIT-1:0] rr_data_132,
        output wire [QNT_BIT-1:0] rr_data_133,
        output wire [QNT_BIT-1:0] rr_data_134,
        output wire [QNT_BIT-1:0] rr_data_135,
        output wire [QNT_BIT-1:0] rr_data_136,
        output wire [QNT_BIT-1:0] rr_data_137,
        output wire [QNT_BIT-1:0] rr_data_138,
        output wire [QNT_BIT-1:0] rr_data_139,
        output wire [QNT_BIT-1:0] rr_data_140,
        output wire [QNT_BIT-1:0] rr_data_141,
        output wire [QNT_BIT-1:0] rr_data_142,
        output wire [QNT_BIT-1:0] rr_data_143,
        output wire [QNT_BIT-1:0] rr_data_144,
        output wire [QNT_BIT-1:0] rr_data_145,
        output wire [QNT_BIT-1:0] rr_data_146,
        output wire [QNT_BIT-1:0] rr_data_147,
        output wire [QNT_BIT-1:0] rr_data_148,
        output wire [QNT_BIT-1:0] rr_data_149,
        output wire [QNT_BIT-1:0] rr_data_150,
        output wire [QNT_BIT-1:0] rr_data_151,
        output wire [QNT_BIT-1:0] rr_data_152,
        output wire [QNT_BIT-1:0] rr_data_153,
        output wire [QNT_BIT-1:0] rr_data_154,
        output wire [QNT_BIT-1:0] rr_data_155,
        output wire [QNT_BIT-1:0] rr_data_156,
        output wire [QNT_BIT-1:0] rr_data_157,
        output wire [QNT_BIT-1:0] rr_data_158,
        output wire [QNT_BIT-1:0] rr_data_159,
        output wire [QNT_BIT-1:0] rr_data_160,
        output wire [QNT_BIT-1:0] rr_data_161,
        output wire [QNT_BIT-1:0] rr_data_162,
        output wire [QNT_BIT-1:0] rr_data_163,
        output wire [QNT_BIT-1:0] rr_data_164,
        output wire [QNT_BIT-1:0] rr_data_165,
        output wire [QNT_BIT-1:0] rr_data_166,
        output wire [QNT_BIT-1:0] rr_data_167,
        output wire [QNT_BIT-1:0] rr_data_168,
        output wire [QNT_BIT-1:0] rr_data_169,
        output wire [QNT_BIT-1:0] rr_data_170,
        output wire [QNT_BIT-1:0] rr_data_171,
        output wire [QNT_BIT-1:0] rr_data_172,
        output wire [QNT_BIT-1:0] rr_data_173,
        output wire [QNT_BIT-1:0] rr_data_174,
        output wire [QNT_BIT-1:0] rr_data_175,
        output wire [QNT_BIT-1:0] rr_data_176,
        output wire [QNT_BIT-1:0] rr_data_177,
        output wire [QNT_BIT-1:0] rr_data_178,
        output wire [QNT_BIT-1:0] rr_data_179,
        output wire [QNT_BIT-1:0] rr_data_180,
        output wire [QNT_BIT-1:0] rr_data_181,
        output wire [QNT_BIT-1:0] rr_data_182,
        output wire [QNT_BIT-1:0] rr_data_183,
        output wire [QNT_BIT-1:0] rr_data_184,
        output wire [QNT_BIT-1:0] rr_data_185,
        output wire [QNT_BIT-1:0] rr_data_186,
        output wire [QNT_BIT-1:0] rr_data_187,
        output wire [QNT_BIT-1:0] rr_data_188,
        output wire [QNT_BIT-1:0] rr_data_189,
        output wire [QNT_BIT-1:0] rr_data_190,
        output wire [QNT_BIT-1:0] rr_data_191,
        output wire [QNT_BIT-1:0] rr_data_192,
        output wire [QNT_BIT-1:0] rr_data_193,
        output wire [QNT_BIT-1:0] rr_data_194,
        output wire [QNT_BIT-1:0] rr_data_195,
        output wire [QNT_BIT-1:0] rr_data_196,
        output wire [QNT_BIT-1:0] rr_data_197,
        output wire [QNT_BIT-1:0] rr_data_198,
        output wire [QNT_BIT-1:0] rr_data_199,
        output wire [QNT_BIT-1:0] rr_data_200,
        output wire [QNT_BIT-1:0] rr_data_201,
        output wire [QNT_BIT-1:0] rr_data_202,
        output wire [QNT_BIT-1:0] rr_data_203,
        output wire [QNT_BIT-1:0] rr_data_204,
        output wire [QNT_BIT-1:0] rr_data_205,
        output wire [QNT_BIT-1:0] rr_data_206,
        output wire [QNT_BIT-1:0] rr_data_207,
        output wire [QNT_BIT-1:0] rr_data_208,
        output wire [QNT_BIT-1:0] rr_data_209,
        output wire [QNT_BIT-1:0] rr_data_210,
        output wire [QNT_BIT-1:0] rr_data_211,
        output wire [QNT_BIT-1:0] rr_data_212,
        output wire [QNT_BIT-1:0] rr_data_213,
        output wire [QNT_BIT-1:0] rr_data_214,
        output wire [QNT_BIT-1:0] rr_data_215,
        output wire [QNT_BIT-1:0] rr_data_216,
        output wire [QNT_BIT-1:0] rr_data_217,
        output wire [QNT_BIT-1:0] rr_data_218,
        output wire [QNT_BIT-1:0] rr_data_219,
        output wire [QNT_BIT-1:0] rr_data_220,
        output wire [QNT_BIT-1:0] rr_data_221,
        output wire [QNT_BIT-1:0] rr_data_222,
        output wire [QNT_BIT-1:0] rr_data_223,
        output wire [QNT_BIT-1:0] rr_data_224,
        output wire [QNT_BIT-1:0] rr_data_225,
        output wire [QNT_BIT-1:0] rr_data_226,
        output wire [QNT_BIT-1:0] rr_data_227,
        output wire [QNT_BIT-1:0] rr_data_228,
        output wire [QNT_BIT-1:0] rr_data_229,
        output wire [QNT_BIT-1:0] rr_data_230,
        output wire [QNT_BIT-1:0] rr_data_231,
        output wire [QNT_BIT-1:0] rr_data_232,
        output wire [QNT_BIT-1:0] rr_data_233,
        output wire [QNT_BIT-1:0] rr_data_234,
        output wire [QNT_BIT-1:0] rr_data_235,
        output wire [QNT_BIT-1:0] rr_data_236,
        output wire [QNT_BIT-1:0] rr_data_237,
        output wire [QNT_BIT-1:0] rr_data_238,
        output wire [QNT_BIT-1:0] rr_data_239,
        output wire [QNT_BIT-1:0] rr_data_240,
        output wire [QNT_BIT-1:0] rr_data_241,
        output wire [QNT_BIT-1:0] rr_data_242,
        output wire [QNT_BIT-1:0] rr_data_243,
        output wire [QNT_BIT-1:0] rr_data_244,
        output wire [QNT_BIT-1:0] rr_data_245,
        output wire [QNT_BIT-1:0] rr_data_246,
        output wire [QNT_BIT-1:0] rr_data_247,
        output wire [QNT_BIT-1:0] rr_data_248,
        output wire [QNT_BIT-1:0] rr_data_249,
        output wire [QNT_BIT-1:0] rr_data_250,
        output wire [QNT_BIT-1:0] rr_data_251,
        output wire [QNT_BIT-1:0] rr_data_252,
        output wire [QNT_BIT-1:0] rr_data_253,
        output wire [QNT_BIT-1:0] rr_data_254,
        output wire [QNT_BIT-1:0] rr_data_255,
        output wire [QNT_BIT-1:0] rr_data_256,
        output wire [QNT_BIT-1:0] rr_data_257,
        output wire [QNT_BIT-1:0] rr_data_258,
        output wire [QNT_BIT-1:0] rr_data_259,
        output wire [QNT_BIT-1:0] rr_data_260,
        output wire [QNT_BIT-1:0] rr_data_261,
        output wire [QNT_BIT-1:0] rr_data_262,
        output wire [QNT_BIT-1:0] rr_data_263,
        output wire [QNT_BIT-1:0] rr_data_264,
        output wire [QNT_BIT-1:0] rr_data_265,
        output wire [QNT_BIT-1:0] rr_data_266,
        output wire [QNT_BIT-1:0] rr_data_267,
        output wire [QNT_BIT-1:0] rr_data_268,
        output wire [QNT_BIT-1:0] rr_data_269,
        output wire [QNT_BIT-1:0] rr_data_270,
        output wire [QNT_BIT-1:0] rr_data_271,
        output wire [QNT_BIT-1:0] rr_data_272,
        output wire [QNT_BIT-1:0] rr_data_273,
        output wire [QNT_BIT-1:0] rr_data_274,
        output wire [QNT_BIT-1:0] rr_data_275,
        output wire [QNT_BIT-1:0] rr_data_276,
        output wire [QNT_BIT-1:0] rr_data_277,
        output wire [QNT_BIT-1:0] rr_data_278,
        output wire [QNT_BIT-1:0] rr_data_279,
        output wire [QNT_BIT-1:0] rr_data_280,
        output wire [QNT_BIT-1:0] rr_data_281,
        output wire [QNT_BIT-1:0] rr_data_282,
        output wire [QNT_BIT-1:0] rr_data_283,
        output wire [QNT_BIT-1:0] rr_data_284,
        output wire [QNT_BIT-1:0] rr_data_285,
        output wire [QNT_BIT-1:0] rr_data_286,
        output wire [QNT_BIT-1:0] rr_data_287,
        output wire [QNT_BIT-1:0] rr_data_288,
        output wire [QNT_BIT-1:0] rr_data_289,
        output wire [QNT_BIT-1:0] rr_data_290,
        output wire [QNT_BIT-1:0] rr_data_291,
        output wire [QNT_BIT-1:0] rr_data_292,
        output wire [QNT_BIT-1:0] rr_data_293,
        output wire [QNT_BIT-1:0] rr_data_294,
        output wire [QNT_BIT-1:0] rr_data_295,
        output wire [QNT_BIT-1:0] rr_data_296,
        output wire [QNT_BIT-1:0] rr_data_297,
        output wire [QNT_BIT-1:0] rr_data_298,
        output wire [QNT_BIT-1:0] rr_data_299,
        output wire [QNT_BIT-1:0] rr_data_300,
        output wire [QNT_BIT-1:0] rr_data_301,
        output wire [QNT_BIT-1:0] rr_data_302,
        output wire [QNT_BIT-1:0] rr_data_303,
        output wire [QNT_BIT-1:0] rr_data_304,
        output wire [QNT_BIT-1:0] rr_data_305,
        output wire [QNT_BIT-1:0] rr_data_306,
        output wire [QNT_BIT-1:0] rr_data_307,
        output wire [QNT_BIT-1:0] rr_data_308,
        output wire [QNT_BIT-1:0] rr_data_309,
        output wire [QNT_BIT-1:0] rr_data_310,
        output wire [QNT_BIT-1:0] rr_data_311,
        output wire [QNT_BIT-1:0] rr_data_312,
        output wire [QNT_BIT-1:0] rr_data_313,
        output wire [QNT_BIT-1:0] rr_data_314,
        output wire [QNT_BIT-1:0] rr_data_315,
        output wire [QNT_BIT-1:0] rr_data_316,
        output wire [QNT_BIT-1:0] rr_data_317,
        output wire [QNT_BIT-1:0] rr_data_318,
        output wire [QNT_BIT-1:0] rr_data_319,
        output wire [QNT_BIT-1:0] rr_data_320,
        output wire [QNT_BIT-1:0] rr_data_321,
        output wire [QNT_BIT-1:0] rr_data_322,
        output wire [QNT_BIT-1:0] rr_data_323,
        output wire [QNT_BIT-1:0] rr_data_324,
        output wire [QNT_BIT-1:0] rr_data_325,
        output wire [QNT_BIT-1:0] rr_data_326,
        output wire [QNT_BIT-1:0] rr_data_327,
        output wire [QNT_BIT-1:0] rr_data_328,
        output wire [QNT_BIT-1:0] rr_data_329,
        output wire [QNT_BIT-1:0] rr_data_330,
        output wire [QNT_BIT-1:0] rr_data_331,
        output wire [QNT_BIT-1:0] rr_data_332,
        output wire [QNT_BIT-1:0] rr_data_333,
        output wire [QNT_BIT-1:0] rr_data_334,
        output wire [QNT_BIT-1:0] rr_data_335,
        output wire [QNT_BIT-1:0] rr_data_336,
        output wire [QNT_BIT-1:0] rr_data_337,
        output wire [QNT_BIT-1:0] rr_data_338,
        output wire [QNT_BIT-1:0] rr_data_339,
        output wire [QNT_BIT-1:0] rr_data_340,
        output wire [QNT_BIT-1:0] rr_data_341,
        output wire [QNT_BIT-1:0] rr_data_342,
        output wire [QNT_BIT-1:0] rr_data_343,
        output wire [QNT_BIT-1:0] rr_data_344,
        output wire [QNT_BIT-1:0] rr_data_345,
        output wire [QNT_BIT-1:0] rr_data_346,
        output wire [QNT_BIT-1:0] rr_data_347,
        output wire [QNT_BIT-1:0] rr_data_348,
        output wire [QNT_BIT-1:0] rr_data_349,
        output wire [QNT_BIT-1:0] rr_data_350,
        output wire [QNT_BIT-1:0] rr_data_351,
        output wire [QNT_BIT-1:0] rr_data_352,
        output wire [QNT_BIT-1:0] rr_data_353,
        output wire [QNT_BIT-1:0] rr_data_354,
        output wire [QNT_BIT-1:0] rr_data_355,
        output wire [QNT_BIT-1:0] rr_data_356,
        output wire [QNT_BIT-1:0] rr_data_357,
        output wire [QNT_BIT-1:0] rr_data_358,
        output wire [QNT_BIT-1:0] rr_data_359,
        output wire [QNT_BIT-1:0] rr_data_360,
        output wire [QNT_BIT-1:0] rr_data_361,
        output wire [QNT_BIT-1:0] rr_data_362,
        output wire [QNT_BIT-1:0] rr_data_363,
        output wire [QNT_BIT-1:0] rr_data_364,
        output wire [QNT_BIT-1:0] rr_data_365,
        output wire [QNT_BIT-1:0] rr_data_366,
        output wire [QNT_BIT-1:0] rr_data_367,
        output wire [QNT_BIT-1:0] rr_data_368,
        output wire [QNT_BIT-1:0] rr_data_369,
        output wire [QNT_BIT-1:0] rr_data_370,
        output wire [QNT_BIT-1:0] rr_data_371,
        output wire [QNT_BIT-1:0] rr_data_372,
        output wire [QNT_BIT-1:0] rr_data_373,
        output wire [QNT_BIT-1:0] rr_data_374,
        output wire [QNT_BIT-1:0] rr_data_375,
        output wire [QNT_BIT-1:0] rr_data_376,
        output wire [QNT_BIT-1:0] rr_data_377,
        output wire [QNT_BIT-1:0] rr_data_378,
        output wire [QNT_BIT-1:0] rr_data_379,
        output wire [QNT_BIT-1:0] rr_data_380,
        output wire [QNT_BIT-1:0] rr_data_381,
        output wire [QNT_BIT-1:0] rr_data_382,
        output wire [QNT_BIT-1:0] rr_data_383,
        output wire [QNT_BIT-1:0] rr_data_384,
        output wire [QNT_BIT-1:0] rr_data_385,
        output wire [QNT_BIT-1:0] rr_data_386,
        output wire [QNT_BIT-1:0] rr_data_387,
        output wire [QNT_BIT-1:0] rr_data_388,
        output wire [QNT_BIT-1:0] rr_data_389,
        output wire [QNT_BIT-1:0] rr_data_390,
        output wire [QNT_BIT-1:0] rr_data_391,
        output wire [QNT_BIT-1:0] rr_data_392,
        output wire [QNT_BIT-1:0] rr_data_393,
        output wire [QNT_BIT-1:0] rr_data_394,
        output wire [QNT_BIT-1:0] rr_data_395,
        output wire [QNT_BIT-1:0] rr_data_396,
        output wire [QNT_BIT-1:0] rr_data_397,
        output wire [QNT_BIT-1:0] rr_data_398,
        output wire [QNT_BIT-1:0] rr_data_399,
        output wire [QNT_BIT-1:0] rr_data_400,
        output wire [QNT_BIT-1:0] rr_data_401,
        output wire [QNT_BIT-1:0] rr_data_402,
        output wire [QNT_BIT-1:0] rr_data_403,
        output wire [QNT_BIT-1:0] rr_data_404,
        output wire [QNT_BIT-1:0] rr_data_405,
        output wire [QNT_BIT-1:0] rr_data_406,
        output wire [QNT_BIT-1:0] rr_data_407,
        output wire [QNT_BIT-1:0] rr_data_408,
        output wire [QNT_BIT-1:0] rr_data_409,
        output wire [QNT_BIT-1:0] rr_data_410,
        output wire [QNT_BIT-1:0] rr_data_411,
        output wire [QNT_BIT-1:0] rr_data_412,
        output wire [QNT_BIT-1:0] rr_data_413,
        output wire [QNT_BIT-1:0] rr_data_414,
        output wire [QNT_BIT-1:0] rr_data_415,
        output wire [QNT_BIT-1:0] rr_data_416,
        output wire [QNT_BIT-1:0] rr_data_417,
        output wire [QNT_BIT-1:0] rr_data_418,
        output wire [QNT_BIT-1:0] rr_data_419,
        output wire [QNT_BIT-1:0] rr_data_420,
        output wire [QNT_BIT-1:0] rr_data_421,
        output wire [QNT_BIT-1:0] rr_data_422,
        output wire [QNT_BIT-1:0] rr_data_423,
        output wire [QNT_BIT-1:0] rr_data_424,
        output wire [QNT_BIT-1:0] rr_data_425,
        output wire [QNT_BIT-1:0] rr_data_426,
        output wire [QNT_BIT-1:0] rr_data_427,
        output wire [QNT_BIT-1:0] rr_data_428,
        output wire [QNT_BIT-1:0] rr_data_429,
        output wire [QNT_BIT-1:0] rr_data_430,
        output wire [QNT_BIT-1:0] rr_data_431,
        output wire [QNT_BIT-1:0] rr_data_432,
        output wire [QNT_BIT-1:0] rr_data_433,
        output wire [QNT_BIT-1:0] rr_data_434,
        output wire [QNT_BIT-1:0] rr_data_435,
        output wire [QNT_BIT-1:0] rr_data_436,
        output wire [QNT_BIT-1:0] rr_data_437,
        output wire [QNT_BIT-1:0] rr_data_438,
        output wire [QNT_BIT-1:0] rr_data_439,
        output wire [QNT_BIT-1:0] rr_data_440,
        output wire [QNT_BIT-1:0] rr_data_441,
        output wire [QNT_BIT-1:0] rr_data_442,
        output wire [QNT_BIT-1:0] rr_data_443,
        output wire [QNT_BIT-1:0] rr_data_444,
        output wire [QNT_BIT-1:0] rr_data_445,
        output wire [QNT_BIT-1:0] rr_data_446,
        output wire [QNT_BIT-1:0] rr_data_447,
        output wire [QNT_BIT-1:0] rr_data_448,
        output wire [QNT_BIT-1:0] rr_data_449,
        output wire [QNT_BIT-1:0] rr_data_450,
        output wire [QNT_BIT-1:0] rr_data_451,
        output wire [QNT_BIT-1:0] rr_data_452,
        output wire [QNT_BIT-1:0] rr_data_453,
        output wire [QNT_BIT-1:0] rr_data_454,
        output wire [QNT_BIT-1:0] rr_data_455,
        output wire [QNT_BIT-1:0] rr_data_456,
        output wire [QNT_BIT-1:0] rr_data_457,
        output wire [QNT_BIT-1:0] rr_data_458,
        output wire [QNT_BIT-1:0] rr_data_459,
        output wire [QNT_BIT-1:0] rr_data_460,
        output wire [QNT_BIT-1:0] rr_data_461,
        output wire [QNT_BIT-1:0] rr_data_462,
        output wire [QNT_BIT-1:0] rr_data_463,
        output wire [QNT_BIT-1:0] rr_data_464,
        output wire [QNT_BIT-1:0] rr_data_465,
        output wire [QNT_BIT-1:0] rr_data_466,
        output wire [QNT_BIT-1:0] rr_data_467,
        output wire [QNT_BIT-1:0] rr_data_468,
        output wire [QNT_BIT-1:0] rr_data_469,
        output wire [QNT_BIT-1:0] rr_data_470,
        output wire [QNT_BIT-1:0] rr_data_471,
        output wire [QNT_BIT-1:0] rr_data_472,
        output wire [QNT_BIT-1:0] rr_data_473,
        output wire [QNT_BIT-1:0] rr_data_474,
        output wire [QNT_BIT-1:0] rr_data_475,
        output wire [QNT_BIT-1:0] rr_data_476,
        output wire [QNT_BIT-1:0] rr_data_477,
        output wire [QNT_BIT-1:0] rr_data_478,
        output wire [QNT_BIT-1:0] rr_data_479,
        output wire [QNT_BIT-1:0] rr_data_480,
        output wire [QNT_BIT-1:0] rr_data_481,
        output wire [QNT_BIT-1:0] rr_data_482,
        output wire [QNT_BIT-1:0] rr_data_483,
        output wire [QNT_BIT-1:0] rr_data_484,
        output wire [QNT_BIT-1:0] rr_data_485,
        output wire [QNT_BIT-1:0] rr_data_486,
        output wire [QNT_BIT-1:0] rr_data_487,
        output wire [QNT_BIT-1:0] rr_data_488,
        output wire [QNT_BIT-1:0] rr_data_489,
        output wire [QNT_BIT-1:0] rr_data_490,
        output wire [QNT_BIT-1:0] rr_data_491,
        output wire [QNT_BIT-1:0] rr_data_492,
        output wire [QNT_BIT-1:0] rr_data_493,
        output wire [QNT_BIT-1:0] rr_data_494,
        output wire [QNT_BIT-1:0] rr_data_495,
        output wire [QNT_BIT-1:0] rr_data_496,
        output wire [QNT_BIT-1:0] rr_data_497,
        output wire [QNT_BIT-1:0] rr_data_498,
        output wire [QNT_BIT-1:0] rr_data_499,
        output wire [QNT_BIT-1:0] rr_data_500,
        output wire [QNT_BIT-1:0] rr_data_501,
        output wire [QNT_BIT-1:0] rr_data_502,
        output wire [QNT_BIT-1:0] rr_data_503,
        output wire [QNT_BIT-1:0] rr_data_504,
        output wire [QNT_BIT-1:0] rr_data_505,
        output wire [QNT_BIT-1:0] rr_data_506,
        output wire [QNT_BIT-1:0] rr_data_507,
        output wire [QNT_BIT-1:0] rr_data_508,
        output wire [QNT_BIT-1:0] rr_data_509,
        output wire [QNT_BIT-1:0] rr_data_510,
        output wire [QNT_BIT-1:0] rr_data_511,
        output wire [QNT_BIT-1:0] rr_data_512,
        output wire [QNT_BIT-1:0] rr_data_513,
        output wire [QNT_BIT-1:0] rr_data_514,
        output wire [QNT_BIT-1:0] rr_data_515,
        output wire [QNT_BIT-1:0] rr_data_516,
        output wire [QNT_BIT-1:0] rr_data_517,
        output wire [QNT_BIT-1:0] rr_data_518,
        output wire [QNT_BIT-1:0] rr_data_519,
        output wire [QNT_BIT-1:0] rr_data_520,
        output wire [QNT_BIT-1:0] rr_data_521,
        output wire [QNT_BIT-1:0] rr_data_522,
        output wire [QNT_BIT-1:0] rr_data_523,
        output wire [QNT_BIT-1:0] rr_data_524,
        output wire [QNT_BIT-1:0] rr_data_525,
        output wire [QNT_BIT-1:0] rr_data_526,
        output wire [QNT_BIT-1:0] rr_data_527,
        output wire [QNT_BIT-1:0] rr_data_528,
        output wire [QNT_BIT-1:0] rr_data_529,
        output wire [QNT_BIT-1:0] rr_data_530,
        output wire [QNT_BIT-1:0] rr_data_531,
        output wire [QNT_BIT-1:0] rr_data_532,
        output wire [QNT_BIT-1:0] rr_data_533

    );

    // * 乒乓操作的存储模块

    reg [QNT_BIT-1:0] page_0[QC_LDPC_COL_COUNT-1:0][QC_LDPC_BLOCK_SIZE-1:0];  // 第 i 个扩展矩阵的第 j 个值
    reg [QNT_BIT-1:0] page_1[QC_LDPC_COL_COUNT-1:0][QC_LDPC_BLOCK_SIZE-1:0];  // 第 i 个扩展矩阵的第 j 个值

    // 初始化与写入逻辑
    integer i, j;
    always @(posedge sys_clk or negedge sys_rst_n) begin
        if (sys_rst_n == 1'b0) begin
            for (i = 0; i < QC_LDPC_COL_COUNT; i = i + 1) begin
                for (j = 0; j < QC_LDPC_BLOCK_SIZE; j = j + 1) begin
                    page_0[i][j] <= {QNT_BIT{1'b0}};
                    page_1[i][j] <= {QNT_BIT{1'b0}};
                end
            end
        end
        else if (write_en) begin
            if (write_page == 1'b0)
                page_0[write_col_cnt][write_cnt] <= sink;
            else
                page_1[write_col_cnt][write_cnt] <= sink;
        end
    end

    genvar i;
    generate
    for (i=1; i<=QC_LDPC_COL_COUNT; i=i+1) begin
        assign rr_data_i = read_page ? page_1[i-1][read_cnt] : page_0[i-1][read_cnt];
    end
    endgenerate











endmodule
