module judge_ctrl (
        input wire sys_clk,
        input wire sys_rst_n,
        input wire flag_judge_start, // ? 控制信号给的

    input wire [63:0] bit_data_1,   // 后验概率的符号位，也就是硬判决的输入
    input wire [63:0] bit_data_2,
    input wire [63:0] bit_data_3,
    input wire [63:0] bit_data_4,
    input wire [63:0] bit_data_5,
    input wire [63:0] bit_data_6,
    input wire [63:0] bit_data_7,
    input wire [63:0] bit_data_8,
    input wire [63:0] bit_data_9,
    input wire [63:0] bit_data_10,
    input wire [63:0] bit_data_11,
    input wire [63:0] bit_data_12,
    input wire [63:0] bit_data_13,
    input wire [63:0] bit_data_14,
    input wire [63:0] bit_data_15,
    input wire [63:0] bit_data_16,
    input wire [63:0] bit_data_17,
    input wire [63:0] bit_data_18,
    input wire [63:0] bit_data_19,
    input wire [63:0] bit_data_20,
    input wire [63:0] bit_data_21,
    input wire [63:0] bit_data_22,
    input wire [63:0] bit_data_23,
    input wire [63:0] bit_data_24,
    input wire [63:0] bit_data_25,
    input wire [63:0] bit_data_26,
    input wire [63:0] bit_data_27,
    input wire [63:0] bit_data_28,
    input wire [63:0] bit_data_29,
    input wire [63:0] bit_data_30,
    input wire [63:0] bit_data_31,
    input wire [63:0] bit_data_32,
    input wire [63:0] bit_data_33,
    input wire [63:0] bit_data_34,
    input wire [63:0] bit_data_35,
    input wire [63:0] bit_data_36,
    input wire [63:0] bit_data_37,
    input wire [63:0] bit_data_38,
    input wire [63:0] bit_data_39,
    input wire [63:0] bit_data_40,
    input wire [63:0] bit_data_41,
    input wire [63:0] bit_data_42,
    input wire [63:0] bit_data_43,
    input wire [63:0] bit_data_44,
    input wire [63:0] bit_data_45,
    input wire [63:0] bit_data_46,
    input wire [63:0] bit_data_47,
    input wire [63:0] bit_data_48,
    input wire [63:0] bit_data_49,
    input wire [63:0] bit_data_50,
    input wire [63:0] bit_data_51,
    input wire [63:0] bit_data_52,
    input wire [63:0] bit_data_53,
    input wire [63:0] bit_data_54,
    input wire [63:0] bit_data_55,
    input wire [63:0] bit_data_56,
    input wire [63:0] bit_data_57,
    input wire [63:0] bit_data_58,
    input wire [63:0] bit_data_59,
    input wire [63:0] bit_data_60,
    input wire [63:0] bit_data_61,
    input wire [63:0] bit_data_62,
    input wire [63:0] bit_data_63,
    input wire [63:0] bit_data_64,
    input wire [63:0] bit_data_65,
    input wire [63:0] bit_data_66,
    input wire [63:0] bit_data_67,
    input wire [63:0] bit_data_68,
    input wire [63:0] bit_data_69,
    input wire [63:0] bit_data_70,
    input wire [63:0] bit_data_71,
    input wire [63:0] bit_data_72,
    input wire [63:0] bit_data_73,
    input wire [63:0] bit_data_74,
    input wire [63:0] bit_data_75,
    input wire [63:0] bit_data_76,
    input wire [63:0] bit_data_77,
    input wire [63:0] bit_data_78,
    input wire [63:0] bit_data_79,
    input wire [63:0] bit_data_80,
    input wire [63:0] bit_data_81,
    input wire [63:0] bit_data_82,
    input wire [63:0] bit_data_83,
    input wire [63:0] bit_data_84,
    input wire [63:0] bit_data_85,
    input wire [63:0] bit_data_86,
    input wire [63:0] bit_data_87,
    input wire [63:0] bit_data_88,
    input wire [63:0] bit_data_89,
    input wire [63:0] bit_data_90,
    input wire [63:0] bit_data_91,
    input wire [63:0] bit_data_92,
    input wire [63:0] bit_data_93,
    input wire [63:0] bit_data_94,
    input wire [63:0] bit_data_95,
    input wire [63:0] bit_data_96,
    input wire [63:0] bit_data_97,
    input wire [63:0] bit_data_98,
    input wire [63:0] bit_data_99,
    input wire [63:0] bit_data_100,
    input wire [63:0] bit_data_101,
    input wire [63:0] bit_data_102,
    input wire [63:0] bit_data_103,
    input wire [63:0] bit_data_104,
    input wire [63:0] bit_data_105,
    input wire [63:0] bit_data_106,
    input wire [63:0] bit_data_107,
    input wire [63:0] bit_data_108,
    input wire [63:0] bit_data_109,
    input wire [63:0] bit_data_110,
    input wire [63:0] bit_data_111,
    input wire [63:0] bit_data_112,
    input wire [63:0] bit_data_113,
    input wire [63:0] bit_data_114,
    input wire [63:0] bit_data_115,
    input wire [63:0] bit_data_116,
    input wire [63:0] bit_data_117,
    input wire [63:0] bit_data_118,
    input wire [63:0] bit_data_119,
    input wire [63:0] bit_data_120,
    input wire [63:0] bit_data_121,
    input wire [63:0] bit_data_122,
    input wire [63:0] bit_data_123,
    input wire [63:0] bit_data_124,
    input wire [63:0] bit_data_125,
    input wire [63:0] bit_data_126,
    input wire [63:0] bit_data_127,
    input wire [63:0] bit_data_128,
    input wire [63:0] bit_data_129,
    input wire [63:0] bit_data_130,
    input wire [63:0] bit_data_131,
    input wire [63:0] bit_data_132,
    input wire [63:0] bit_data_133,
    input wire [63:0] bit_data_134,
    input wire [63:0] bit_data_135,
    input wire [63:0] bit_data_136,
    input wire [63:0] bit_data_137,
    input wire [63:0] bit_data_138,
    input wire [63:0] bit_data_139,
    input wire [63:0] bit_data_140,
    input wire [63:0] bit_data_141,
    input wire [63:0] bit_data_142,
    input wire [63:0] bit_data_143,
    input wire [63:0] bit_data_144,
    input wire [63:0] bit_data_145,
    input wire [63:0] bit_data_146,
    input wire [63:0] bit_data_147,
    input wire [63:0] bit_data_148,
    input wire [63:0] bit_data_149,
    input wire [63:0] bit_data_150,
    input wire [63:0] bit_data_151,
    input wire [63:0] bit_data_152,
    input wire [63:0] bit_data_153,
    input wire [63:0] bit_data_154,
    input wire [63:0] bit_data_155,
    input wire [63:0] bit_data_156,
    input wire [63:0] bit_data_157,
    input wire [63:0] bit_data_158,
    input wire [63:0] bit_data_159,
    input wire [63:0] bit_data_160,
    input wire [63:0] bit_data_161,
    input wire [63:0] bit_data_162,
    input wire [63:0] bit_data_163,
    input wire [63:0] bit_data_164,
    input wire [63:0] bit_data_165,
    input wire [63:0] bit_data_166,
    input wire [63:0] bit_data_167,
    input wire [63:0] bit_data_168,
    input wire [63:0] bit_data_169,
    input wire [63:0] bit_data_170,
    input wire [63:0] bit_data_171,
    input wire [63:0] bit_data_172,
    input wire [63:0] bit_data_173,
    input wire [63:0] bit_data_174,
    input wire [63:0] bit_data_175,
    input wire [63:0] bit_data_176,
    input wire [63:0] bit_data_177,
    input wire [63:0] bit_data_178,
    input wire [63:0] bit_data_179,
    input wire [63:0] bit_data_180,
    input wire [63:0] bit_data_181,
    input wire [63:0] bit_data_182,
    input wire [63:0] bit_data_183,
    input wire [63:0] bit_data_184,
    input wire [63:0] bit_data_185,
    input wire [63:0] bit_data_186,
    input wire [63:0] bit_data_187,
    input wire [63:0] bit_data_188,
    input wire [63:0] bit_data_189,
    input wire [63:0] bit_data_190,
    input wire [63:0] bit_data_191,
    input wire [63:0] bit_data_192,
    input wire [63:0] bit_data_193,
    input wire [63:0] bit_data_194,
    input wire [63:0] bit_data_195,
    input wire [63:0] bit_data_196,
    input wire [63:0] bit_data_197,
    input wire [63:0] bit_data_198,
    input wire [63:0] bit_data_199,
    input wire [63:0] bit_data_200,
    input wire [63:0] bit_data_201,
    input wire [63:0] bit_data_202,
    input wire [63:0] bit_data_203,
    input wire [63:0] bit_data_204,
    input wire [63:0] bit_data_205,
    input wire [63:0] bit_data_206,
    input wire [63:0] bit_data_207,
    input wire [63:0] bit_data_208,
    input wire [63:0] bit_data_209,
    input wire [63:0] bit_data_210,
    input wire [63:0] bit_data_211,
    input wire [63:0] bit_data_212,
    input wire [63:0] bit_data_213,
    input wire [63:0] bit_data_214,
    input wire [63:0] bit_data_215,
    input wire [63:0] bit_data_216,
    input wire [63:0] bit_data_217,
    input wire [63:0] bit_data_218,
    input wire [63:0] bit_data_219,
    input wire [63:0] bit_data_220,
    input wire [63:0] bit_data_221,
    input wire [63:0] bit_data_222,
    input wire [63:0] bit_data_223,
    input wire [63:0] bit_data_224,
    input wire [63:0] bit_data_225,
    input wire [63:0] bit_data_226,
    input wire [63:0] bit_data_227,
    input wire [63:0] bit_data_228,
    input wire [63:0] bit_data_229,
    input wire [63:0] bit_data_230,
    input wire [63:0] bit_data_231,
    input wire [63:0] bit_data_232,
    input wire [63:0] bit_data_233,
    input wire [63:0] bit_data_234,
    input wire [63:0] bit_data_235,
    input wire [63:0] bit_data_236,
    input wire [63:0] bit_data_237,
    input wire [63:0] bit_data_238,
    input wire [63:0] bit_data_239,
    input wire [63:0] bit_data_240,
    input wire [63:0] bit_data_241,
    input wire [63:0] bit_data_242,
    input wire [63:0] bit_data_243,
    input wire [63:0] bit_data_244,
    input wire [63:0] bit_data_245,
    input wire [63:0] bit_data_246,
    input wire [63:0] bit_data_247,
    input wire [63:0] bit_data_248,
    input wire [63:0] bit_data_249,
    input wire [63:0] bit_data_250,
    input wire [63:0] bit_data_251,
    input wire [63:0] bit_data_252,
    input wire [63:0] bit_data_253,
    input wire [63:0] bit_data_254,
    input wire [63:0] bit_data_255,
    input wire [63:0] bit_data_256,
    input wire [63:0] bit_data_257,
    input wire [63:0] bit_data_258,
    input wire [63:0] bit_data_259,
    input wire [63:0] bit_data_260,
    input wire [63:0] bit_data_261,
    input wire [63:0] bit_data_262,
    input wire [63:0] bit_data_263,
    input wire [63:0] bit_data_264,
    input wire [63:0] bit_data_265,
    input wire [63:0] bit_data_266,
    input wire [63:0] bit_data_267,
    input wire [63:0] bit_data_268,
    input wire [63:0] bit_data_269,
    input wire [63:0] bit_data_270,
    input wire [63:0] bit_data_271,
    input wire [63:0] bit_data_272,
    input wire [63:0] bit_data_273,
    input wire [63:0] bit_data_274,
    input wire [63:0] bit_data_275,
    input wire [63:0] bit_data_276,
    input wire [63:0] bit_data_277,
    input wire [63:0] bit_data_278,
    input wire [63:0] bit_data_279,
    input wire [63:0] bit_data_280,
    input wire [63:0] bit_data_281,
    input wire [63:0] bit_data_282,
    input wire [63:0] bit_data_283,
    input wire [63:0] bit_data_284,
    input wire [63:0] bit_data_285,
    input wire [63:0] bit_data_286,
    input wire [63:0] bit_data_287,
    input wire [63:0] bit_data_288,
    input wire [63:0] bit_data_289,
    input wire [63:0] bit_data_290,
    input wire [63:0] bit_data_291,
    input wire [63:0] bit_data_292,
    input wire [63:0] bit_data_293,
    input wire [63:0] bit_data_294,
    input wire [63:0] bit_data_295,
    input wire [63:0] bit_data_296,
    input wire [63:0] bit_data_297,
    input wire [63:0] bit_data_298,
    input wire [63:0] bit_data_299,
    input wire [63:0] bit_data_300,
    input wire [63:0] bit_data_301,
    input wire [63:0] bit_data_302,
    input wire [63:0] bit_data_303,
    input wire [63:0] bit_data_304,
    input wire [63:0] bit_data_305,
    input wire [63:0] bit_data_306,
    input wire [63:0] bit_data_307,
    input wire [63:0] bit_data_308,
    input wire [63:0] bit_data_309,
    input wire [63:0] bit_data_310,
    input wire [63:0] bit_data_311,
    input wire [63:0] bit_data_312,
    input wire [63:0] bit_data_313,
    input wire [63:0] bit_data_314,
    input wire [63:0] bit_data_315,
    input wire [63:0] bit_data_316,
    input wire [63:0] bit_data_317,
    input wire [63:0] bit_data_318,
    input wire [63:0] bit_data_319,
    input wire [63:0] bit_data_320,
    input wire [63:0] bit_data_321,
    input wire [63:0] bit_data_322,
    input wire [63:0] bit_data_323,
    input wire [63:0] bit_data_324,
    input wire [63:0] bit_data_325,
    input wire [63:0] bit_data_326,
    input wire [63:0] bit_data_327,
    input wire [63:0] bit_data_328,
    input wire [63:0] bit_data_329,
    input wire [63:0] bit_data_330,
    input wire [63:0] bit_data_331,
    input wire [63:0] bit_data_332,
    input wire [63:0] bit_data_333,
    input wire [63:0] bit_data_334,
    input wire [63:0] bit_data_335,
    input wire [63:0] bit_data_336,
    input wire [63:0] bit_data_337,
    input wire [63:0] bit_data_338,
    input wire [63:0] bit_data_339,
    input wire [63:0] bit_data_340,
    input wire [63:0] bit_data_341,
    input wire [63:0] bit_data_342,
    input wire [63:0] bit_data_343,
    input wire [63:0] bit_data_344,
    input wire [63:0] bit_data_345,
    input wire [63:0] bit_data_346,
    input wire [63:0] bit_data_347,
    input wire [63:0] bit_data_348,
    input wire [63:0] bit_data_349,
    input wire [63:0] bit_data_350,
    input wire [63:0] bit_data_351,
    input wire [63:0] bit_data_352,
    input wire [63:0] bit_data_353,
    input wire [63:0] bit_data_354,
    input wire [63:0] bit_data_355,
    input wire [63:0] bit_data_356,
    input wire [63:0] bit_data_357,
    input wire [63:0] bit_data_358,
    input wire [63:0] bit_data_359,
    input wire [63:0] bit_data_360,
    input wire [63:0] bit_data_361,
    input wire [63:0] bit_data_362,
    input wire [63:0] bit_data_363,
    input wire [63:0] bit_data_364,
    input wire [63:0] bit_data_365,
    input wire [63:0] bit_data_366,
    input wire [63:0] bit_data_367,
    input wire [63:0] bit_data_368,
    input wire [63:0] bit_data_369,
    input wire [63:0] bit_data_370,
    input wire [63:0] bit_data_371,
    input wire [63:0] bit_data_372,
    input wire [63:0] bit_data_373,
    input wire [63:0] bit_data_374,
    input wire [63:0] bit_data_375,
    input wire [63:0] bit_data_376,
    input wire [63:0] bit_data_377,
    input wire [63:0] bit_data_378,
    input wire [63:0] bit_data_379,
    input wire [63:0] bit_data_380,
    input wire [63:0] bit_data_381,
    input wire [63:0] bit_data_382,
    input wire [63:0] bit_data_383,
    input wire [63:0] bit_data_384,
    input wire [63:0] bit_data_385,
    input wire [63:0] bit_data_386,
    input wire [63:0] bit_data_387,
    input wire [63:0] bit_data_388,
    input wire [63:0] bit_data_389,
    input wire [63:0] bit_data_390,
    input wire [63:0] bit_data_391,
    input wire [63:0] bit_data_392,
    input wire [63:0] bit_data_393,
    input wire [63:0] bit_data_394,
    input wire [63:0] bit_data_395,
    input wire [63:0] bit_data_396,
    input wire [63:0] bit_data_397,
    input wire [63:0] bit_data_398,
    input wire [63:0] bit_data_399,
    input wire [63:0] bit_data_400,
    input wire [63:0] bit_data_401,
    input wire [63:0] bit_data_402,
    input wire [63:0] bit_data_403,
    input wire [63:0] bit_data_404,
    input wire [63:0] bit_data_405,
    input wire [63:0] bit_data_406,
    input wire [63:0] bit_data_407,
    input wire [63:0] bit_data_408,
    input wire [63:0] bit_data_409,
    input wire [63:0] bit_data_410,
    input wire [63:0] bit_data_411,
    input wire [63:0] bit_data_412,
    input wire [63:0] bit_data_413,
    input wire [63:0] bit_data_414,
    input wire [63:0] bit_data_415,
    input wire [63:0] bit_data_416,
    input wire [63:0] bit_data_417,
    input wire [63:0] bit_data_418,
    input wire [63:0] bit_data_419,
    input wire [63:0] bit_data_420,
    input wire [63:0] bit_data_421,
    input wire [63:0] bit_data_422,
    input wire [63:0] bit_data_423,
    input wire [63:0] bit_data_424,
    input wire [63:0] bit_data_425,
    input wire [63:0] bit_data_426,
    input wire [63:0] bit_data_427,
    input wire [63:0] bit_data_428,
    input wire [63:0] bit_data_429,
    input wire [63:0] bit_data_430,
    input wire [63:0] bit_data_431,
    input wire [63:0] bit_data_432,
    input wire [63:0] bit_data_433,
    input wire [63:0] bit_data_434,
    input wire [63:0] bit_data_435,
    input wire [63:0] bit_data_436,
    input wire [63:0] bit_data_437,
    input wire [63:0] bit_data_438,
    input wire [63:0] bit_data_439,
    input wire [63:0] bit_data_440,
    input wire [63:0] bit_data_441,
    input wire [63:0] bit_data_442,
    input wire [63:0] bit_data_443,
    input wire [63:0] bit_data_444,
    input wire [63:0] bit_data_445,
    input wire [63:0] bit_data_446,
    input wire [63:0] bit_data_447,
    input wire [63:0] bit_data_448,
    input wire [63:0] bit_data_449,
    input wire [63:0] bit_data_450,
    input wire [63:0] bit_data_451,
    input wire [63:0] bit_data_452,
    input wire [63:0] bit_data_453,
    input wire [63:0] bit_data_454,
    input wire [63:0] bit_data_455,
    input wire [63:0] bit_data_456,
    input wire [63:0] bit_data_457,
    input wire [63:0] bit_data_458,
    input wire [63:0] bit_data_459,
    input wire [63:0] bit_data_460,
    input wire [63:0] bit_data_461,
    input wire [63:0] bit_data_462,
    input wire [63:0] bit_data_463,
    input wire [63:0] bit_data_464,
    input wire [63:0] bit_data_465,
    input wire [63:0] bit_data_466,
    input wire [63:0] bit_data_467,
    input wire [63:0] bit_data_468,
    input wire [63:0] bit_data_469,
    input wire [63:0] bit_data_470,
    input wire [63:0] bit_data_471,
    input wire [63:0] bit_data_472,
    input wire [63:0] bit_data_473,
    input wire [63:0] bit_data_474,
    input wire [63:0] bit_data_475,
    input wire [63:0] bit_data_476,
    input wire [63:0] bit_data_477,
    input wire [63:0] bit_data_478,
    input wire [63:0] bit_data_479,
    input wire [63:0] bit_data_480,
    input wire [63:0] bit_data_481,
    input wire [63:0] bit_data_482,
    input wire [63:0] bit_data_483,
    input wire [63:0] bit_data_484,
    input wire [63:0] bit_data_485,
    input wire [63:0] bit_data_486,
    input wire [63:0] bit_data_487,
    input wire [63:0] bit_data_488,
    input wire [63:0] bit_data_489,
    input wire [63:0] bit_data_490,
    input wire [63:0] bit_data_491,
    input wire [63:0] bit_data_492,
    input wire [63:0] bit_data_493,
    input wire [63:0] bit_data_494,
    input wire [63:0] bit_data_495,
    input wire [63:0] bit_data_496,
    input wire [63:0] bit_data_497,
    input wire [63:0] bit_data_498,
    input wire [63:0] bit_data_499,
    input wire [63:0] bit_data_500,
    input wire [63:0] bit_data_501,
    input wire [63:0] bit_data_502,
    input wire [63:0] bit_data_503,
    input wire [63:0] bit_data_504,
    input wire [63:0] bit_data_505,
    input wire [63:0] bit_data_506,
    input wire [63:0] bit_data_507,
    input wire [63:0] bit_data_508,
    input wire [63:0] bit_data_509,
    input wire [63:0] bit_data_510,
    input wire [63:0] bit_data_511,
    input wire [63:0] bit_data_512,
    input wire [63:0] bit_data_513,
    input wire [63:0] bit_data_514,
    input wire [63:0] bit_data_515,
    input wire [63:0] bit_data_516,
    input wire [63:0] bit_data_517,
    input wire [63:0] bit_data_518,
    input wire [63:0] bit_data_519,
    input wire [63:0] bit_data_520,
    input wire [63:0] bit_data_521,
    input wire [63:0] bit_data_522,
    input wire [63:0] bit_data_523,
    input wire [63:0] bit_data_524,
    input wire [63:0] bit_data_525,
    input wire [63:0] bit_data_526,
    input wire [63:0] bit_data_527,
    input wire [63:0] bit_data_528,
    input wire [63:0] bit_data_529,
    input wire [63:0] bit_data_530,
    input wire [63:0] bit_data_531,
    input wire [63:0] bit_data_532,
    input wire [63:0] bit_data_533,

        output reg       flag_judge_end,    //判决模块完成
        output reg [6:0] H_sum
    );

    // * 本模块进行判断硬判决的结果正确性


    // 扩展矩阵
`include "Hb_H_QC_N68224_K65536_R0.96_z128.txt"
    /* parameter  cyclic_shif_data_1_2   =   5'd23; */


    reg        judge_en;
    reg        judge_en_reg;
    reg [ 6:0] cnt;
    reg [20:0] judge_bit;  //判断每个校验方程
    reg [ 6:0] judge_sum;


    // wire 定义
`include "addr_shif_define_4KB.txt"
    /* wire	[5:0]	addr_shif_1_2; */


	// 开始进行 judge 操作
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            judge_en <= 1'b0;
    else if (cnt == 7'd63)
            judge_en <= 1'b0;
        else if (flag_judge_start == 1'b1)
            judge_en <= 1'b1;
        else
            judge_en <= judge_en;


    // 给 judge_en_reg 再打一拍
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            judge_en_reg <= 1'b0;
        else
            judge_en_reg <= judge_en;


    // 判断什么时候终止
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            flag_judge_end <= 1'b0;
        else if (judge_en_reg == 1'b1 && judge_en == 1'b0)
            flag_judge_end <= 1'b1;
        else
            flag_judge_end <= 1'b0;


    // 选择判断数据的地址自增器，一个周期并行校验 12 个在不同循环体的校验方程
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            cnt <= 7'd0;
    else if (flag_judge_start == 1'b1 || cnt == 7'd63)
            cnt <= 7'd0;
        else if (judge_en == 1'b1)
            cnt <= cnt + 1'd1;
        else
            cnt <= cnt;


    // 对不满足的校验方程单位（每 12 个为一个单位）数量进行求和
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            judge_sum <= 4'd0;
        else if (flag_judge_start == 1'b1)
            judge_sum <= 4'd0;
        else if (judge_en == 1'b1)
            judge_sum <= judge_sum + judge_bit[0] + judge_bit[1] + judge_bit[2] + judge_bit[3] + judge_bit[4] + judge_bit[5] + judge_bit[6] + judge_bit[7] + judge_bit[8] + judge_bit[9] + judge_bit[10] + judge_bit[11] + judge_bit[12] + judge_bit[13] + judge_bit[14] + judge_bit[15] + judge_bit[16] + judge_bit[17] + judge_bit[18] + judge_bit[19] + judge_bit[20];
        else
            judge_sum <= judge_sum;


    // 对校验结果进行更新
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            H_sum <= 4'd0;
        else if (judge_en_reg == 1'b1 && judge_en == 1'b0)
            H_sum <= judge_sum;
        else
            H_sum <= H_sum;


    // 校验方程的校验结果，即求和判断是否为 0
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            judge_bit <= 21'd0;
        else if (flag_judge_start == 1'b1)
            judge_bit <= 21'd0;
        else if (judge_en == 1'b1) begin
`include "judge_bit_data_4KB.txt"
            /*judge_bit[0]<=	bit_data_2[addr_shif_1_2]+bit_data_3[addr_shif_1_3]+bit_data_9[addr_shif_1_9]+
                  bit_data_10[addr_shif_1_10]+bit_data_13[addr_shif_1_13]+bit_data_14[addr_shif_1_14]; */
        end
        else
            judge_bit <= judge_bit;


    // 根据校验进程和 H 矩阵的扩展因子，计算的校验参与数据在校验循环体中的地址
`include "addr_shif_data_4KB.txt"
    /* assign	addr_shif_1_2=(judge_en==1'b1)?
    ((cnt+cyclic_shif_data_1_2>=6'd24)?
    (cnt-cyclic+shif_data_1_2-6'd24):
    (cnt+cyclic_shif_data_1_2)):6'd0; */

endmodule
