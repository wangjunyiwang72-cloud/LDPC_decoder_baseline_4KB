module buffer_out #(
    parameter QC_LDPC_COL_COUNT = 533
) (
        input wire sys_clk,
        input wire sys_rst_n,
        input wire flag_serial, // ? 控制信号给的，拉高一个周期说明计算完成

    input wire [63:0] bit_data_1,   // 后验概率的符号位，也就是硬判决的输入
    input wire [63:0] bit_data_2,
    input wire [63:0] bit_data_3,
    input wire [63:0] bit_data_4,
    input wire [63:0] bit_data_5,
    input wire [63:0] bit_data_6,
    input wire [63:0] bit_data_7,
    input wire [63:0] bit_data_8,
    input wire [63:0] bit_data_9,
    input wire [63:0] bit_data_10,
    input wire [63:0] bit_data_11,
    input wire [63:0] bit_data_12,
    input wire [63:0] bit_data_13,
    input wire [63:0] bit_data_14,
    input wire [63:0] bit_data_15,
    input wire [63:0] bit_data_16,
    input wire [63:0] bit_data_17,
    input wire [63:0] bit_data_18,
    input wire [63:0] bit_data_19,
    input wire [63:0] bit_data_20,
    input wire [63:0] bit_data_21,
    input wire [63:0] bit_data_22,
    input wire [63:0] bit_data_23,
    input wire [63:0] bit_data_24,
    input wire [63:0] bit_data_25,
    input wire [63:0] bit_data_26,
    input wire [63:0] bit_data_27,
    input wire [63:0] bit_data_28,
    input wire [63:0] bit_data_29,
    input wire [63:0] bit_data_30,
    input wire [63:0] bit_data_31,
    input wire [63:0] bit_data_32,
    input wire [63:0] bit_data_33,
    input wire [63:0] bit_data_34,
    input wire [63:0] bit_data_35,
    input wire [63:0] bit_data_36,
    input wire [63:0] bit_data_37,
    input wire [63:0] bit_data_38,
    input wire [63:0] bit_data_39,
    input wire [63:0] bit_data_40,
    input wire [63:0] bit_data_41,
    input wire [63:0] bit_data_42,
    input wire [63:0] bit_data_43,
    input wire [63:0] bit_data_44,
    input wire [63:0] bit_data_45,
    input wire [63:0] bit_data_46,
    input wire [63:0] bit_data_47,
    input wire [63:0] bit_data_48,
    input wire [63:0] bit_data_49,
    input wire [63:0] bit_data_50,
    input wire [63:0] bit_data_51,
    input wire [63:0] bit_data_52,
    input wire [63:0] bit_data_53,
    input wire [63:0] bit_data_54,
    input wire [63:0] bit_data_55,
    input wire [63:0] bit_data_56,
    input wire [63:0] bit_data_57,
    input wire [63:0] bit_data_58,
    input wire [63:0] bit_data_59,
    input wire [63:0] bit_data_60,
    input wire [63:0] bit_data_61,
    input wire [63:0] bit_data_62,
    input wire [63:0] bit_data_63,
    input wire [63:0] bit_data_64,
    input wire [63:0] bit_data_65,
    input wire [63:0] bit_data_66,
    input wire [63:0] bit_data_67,
    input wire [63:0] bit_data_68,
    input wire [63:0] bit_data_69,
    input wire [63:0] bit_data_70,
    input wire [63:0] bit_data_71,
    input wire [63:0] bit_data_72,
    input wire [63:0] bit_data_73,
    input wire [63:0] bit_data_74,
    input wire [63:0] bit_data_75,
    input wire [63:0] bit_data_76,
    input wire [63:0] bit_data_77,
    input wire [63:0] bit_data_78,
    input wire [63:0] bit_data_79,
    input wire [63:0] bit_data_80,
    input wire [63:0] bit_data_81,
    input wire [63:0] bit_data_82,
    input wire [63:0] bit_data_83,
    input wire [63:0] bit_data_84,
    input wire [63:0] bit_data_85,
    input wire [63:0] bit_data_86,
    input wire [63:0] bit_data_87,
    input wire [63:0] bit_data_88,
    input wire [63:0] bit_data_89,
    input wire [63:0] bit_data_90,
    input wire [63:0] bit_data_91,
    input wire [63:0] bit_data_92,
    input wire [63:0] bit_data_93,
    input wire [63:0] bit_data_94,
    input wire [63:0] bit_data_95,
    input wire [63:0] bit_data_96,
    input wire [63:0] bit_data_97,
    input wire [63:0] bit_data_98,
    input wire [63:0] bit_data_99,
    input wire [63:0] bit_data_100,
    input wire [63:0] bit_data_101,
    input wire [63:0] bit_data_102,
    input wire [63:0] bit_data_103,
    input wire [63:0] bit_data_104,
    input wire [63:0] bit_data_105,
    input wire [63:0] bit_data_106,
    input wire [63:0] bit_data_107,
    input wire [63:0] bit_data_108,
    input wire [63:0] bit_data_109,
    input wire [63:0] bit_data_110,
    input wire [63:0] bit_data_111,
    input wire [63:0] bit_data_112,
    input wire [63:0] bit_data_113,
    input wire [63:0] bit_data_114,
    input wire [63:0] bit_data_115,
    input wire [63:0] bit_data_116,
    input wire [63:0] bit_data_117,
    input wire [63:0] bit_data_118,
    input wire [63:0] bit_data_119,
    input wire [63:0] bit_data_120,
    input wire [63:0] bit_data_121,
    input wire [63:0] bit_data_122,
    input wire [63:0] bit_data_123,
    input wire [63:0] bit_data_124,
    input wire [63:0] bit_data_125,
    input wire [63:0] bit_data_126,
    input wire [63:0] bit_data_127,
    input wire [63:0] bit_data_128,
    input wire [63:0] bit_data_129,
    input wire [63:0] bit_data_130,
    input wire [63:0] bit_data_131,
    input wire [63:0] bit_data_132,
    input wire [63:0] bit_data_133,
    input wire [63:0] bit_data_134,
    input wire [63:0] bit_data_135,
    input wire [63:0] bit_data_136,
    input wire [63:0] bit_data_137,
    input wire [63:0] bit_data_138,
    input wire [63:0] bit_data_139,
    input wire [63:0] bit_data_140,
    input wire [63:0] bit_data_141,
    input wire [63:0] bit_data_142,
    input wire [63:0] bit_data_143,
    input wire [63:0] bit_data_144,
    input wire [63:0] bit_data_145,
    input wire [63:0] bit_data_146,
    input wire [63:0] bit_data_147,
    input wire [63:0] bit_data_148,
    input wire [63:0] bit_data_149,
    input wire [63:0] bit_data_150,
    input wire [63:0] bit_data_151,
    input wire [63:0] bit_data_152,
    input wire [63:0] bit_data_153,
    input wire [63:0] bit_data_154,
    input wire [63:0] bit_data_155,
    input wire [63:0] bit_data_156,
    input wire [63:0] bit_data_157,
    input wire [63:0] bit_data_158,
    input wire [63:0] bit_data_159,
    input wire [63:0] bit_data_160,
    input wire [63:0] bit_data_161,
    input wire [63:0] bit_data_162,
    input wire [63:0] bit_data_163,
    input wire [63:0] bit_data_164,
    input wire [63:0] bit_data_165,
    input wire [63:0] bit_data_166,
    input wire [63:0] bit_data_167,
    input wire [63:0] bit_data_168,
    input wire [63:0] bit_data_169,
    input wire [63:0] bit_data_170,
    input wire [63:0] bit_data_171,
    input wire [63:0] bit_data_172,
    input wire [63:0] bit_data_173,
    input wire [63:0] bit_data_174,
    input wire [63:0] bit_data_175,
    input wire [63:0] bit_data_176,
    input wire [63:0] bit_data_177,
    input wire [63:0] bit_data_178,
    input wire [63:0] bit_data_179,
    input wire [63:0] bit_data_180,
    input wire [63:0] bit_data_181,
    input wire [63:0] bit_data_182,
    input wire [63:0] bit_data_183,
    input wire [63:0] bit_data_184,
    input wire [63:0] bit_data_185,
    input wire [63:0] bit_data_186,
    input wire [63:0] bit_data_187,
    input wire [63:0] bit_data_188,
    input wire [63:0] bit_data_189,
    input wire [63:0] bit_data_190,
    input wire [63:0] bit_data_191,
    input wire [63:0] bit_data_192,
    input wire [63:0] bit_data_193,
    input wire [63:0] bit_data_194,
    input wire [63:0] bit_data_195,
    input wire [63:0] bit_data_196,
    input wire [63:0] bit_data_197,
    input wire [63:0] bit_data_198,
    input wire [63:0] bit_data_199,
    input wire [63:0] bit_data_200,
    input wire [63:0] bit_data_201,
    input wire [63:0] bit_data_202,
    input wire [63:0] bit_data_203,
    input wire [63:0] bit_data_204,
    input wire [63:0] bit_data_205,
    input wire [63:0] bit_data_206,
    input wire [63:0] bit_data_207,
    input wire [63:0] bit_data_208,
    input wire [63:0] bit_data_209,
    input wire [63:0] bit_data_210,
    input wire [63:0] bit_data_211,
    input wire [63:0] bit_data_212,
    input wire [63:0] bit_data_213,
    input wire [63:0] bit_data_214,
    input wire [63:0] bit_data_215,
    input wire [63:0] bit_data_216,
    input wire [63:0] bit_data_217,
    input wire [63:0] bit_data_218,
    input wire [63:0] bit_data_219,
    input wire [63:0] bit_data_220,
    input wire [63:0] bit_data_221,
    input wire [63:0] bit_data_222,
    input wire [63:0] bit_data_223,
    input wire [63:0] bit_data_224,
    input wire [63:0] bit_data_225,
    input wire [63:0] bit_data_226,
    input wire [63:0] bit_data_227,
    input wire [63:0] bit_data_228,
    input wire [63:0] bit_data_229,
    input wire [63:0] bit_data_230,
    input wire [63:0] bit_data_231,
    input wire [63:0] bit_data_232,
    input wire [63:0] bit_data_233,
    input wire [63:0] bit_data_234,
    input wire [63:0] bit_data_235,
    input wire [63:0] bit_data_236,
    input wire [63:0] bit_data_237,
    input wire [63:0] bit_data_238,
    input wire [63:0] bit_data_239,
    input wire [63:0] bit_data_240,
    input wire [63:0] bit_data_241,
    input wire [63:0] bit_data_242,
    input wire [63:0] bit_data_243,
    input wire [63:0] bit_data_244,
    input wire [63:0] bit_data_245,
    input wire [63:0] bit_data_246,
    input wire [63:0] bit_data_247,
    input wire [63:0] bit_data_248,
    input wire [63:0] bit_data_249,
    input wire [63:0] bit_data_250,
    input wire [63:0] bit_data_251,
    input wire [63:0] bit_data_252,
    input wire [63:0] bit_data_253,
    input wire [63:0] bit_data_254,
    input wire [63:0] bit_data_255,
    input wire [63:0] bit_data_256,
    input wire [63:0] bit_data_257,
    input wire [63:0] bit_data_258,
    input wire [63:0] bit_data_259,
    input wire [63:0] bit_data_260,
    input wire [63:0] bit_data_261,
    input wire [63:0] bit_data_262,
    input wire [63:0] bit_data_263,
    input wire [63:0] bit_data_264,
    input wire [63:0] bit_data_265,
    input wire [63:0] bit_data_266,
    input wire [63:0] bit_data_267,
    input wire [63:0] bit_data_268,
    input wire [63:0] bit_data_269,
    input wire [63:0] bit_data_270,
    input wire [63:0] bit_data_271,
    input wire [63:0] bit_data_272,
    input wire [63:0] bit_data_273,
    input wire [63:0] bit_data_274,
    input wire [63:0] bit_data_275,
    input wire [63:0] bit_data_276,
    input wire [63:0] bit_data_277,
    input wire [63:0] bit_data_278,
    input wire [63:0] bit_data_279,
    input wire [63:0] bit_data_280,
    input wire [63:0] bit_data_281,
    input wire [63:0] bit_data_282,
    input wire [63:0] bit_data_283,
    input wire [63:0] bit_data_284,
    input wire [63:0] bit_data_285,
    input wire [63:0] bit_data_286,
    input wire [63:0] bit_data_287,
    input wire [63:0] bit_data_288,
    input wire [63:0] bit_data_289,
    input wire [63:0] bit_data_290,
    input wire [63:0] bit_data_291,
    input wire [63:0] bit_data_292,
    input wire [63:0] bit_data_293,
    input wire [63:0] bit_data_294,
    input wire [63:0] bit_data_295,
    input wire [63:0] bit_data_296,
    input wire [63:0] bit_data_297,
    input wire [63:0] bit_data_298,
    input wire [63:0] bit_data_299,
    input wire [63:0] bit_data_300,
    input wire [63:0] bit_data_301,
    input wire [63:0] bit_data_302,
    input wire [63:0] bit_data_303,
    input wire [63:0] bit_data_304,
    input wire [63:0] bit_data_305,
    input wire [63:0] bit_data_306,
    input wire [63:0] bit_data_307,
    input wire [63:0] bit_data_308,
    input wire [63:0] bit_data_309,
    input wire [63:0] bit_data_310,
    input wire [63:0] bit_data_311,
    input wire [63:0] bit_data_312,
    input wire [63:0] bit_data_313,
    input wire [63:0] bit_data_314,
    input wire [63:0] bit_data_315,
    input wire [63:0] bit_data_316,
    input wire [63:0] bit_data_317,
    input wire [63:0] bit_data_318,
    input wire [63:0] bit_data_319,
    input wire [63:0] bit_data_320,
    input wire [63:0] bit_data_321,
    input wire [63:0] bit_data_322,
    input wire [63:0] bit_data_323,
    input wire [63:0] bit_data_324,
    input wire [63:0] bit_data_325,
    input wire [63:0] bit_data_326,
    input wire [63:0] bit_data_327,
    input wire [63:0] bit_data_328,
    input wire [63:0] bit_data_329,
    input wire [63:0] bit_data_330,
    input wire [63:0] bit_data_331,
    input wire [63:0] bit_data_332,
    input wire [63:0] bit_data_333,
    input wire [63:0] bit_data_334,
    input wire [63:0] bit_data_335,
    input wire [63:0] bit_data_336,
    input wire [63:0] bit_data_337,
    input wire [63:0] bit_data_338,
    input wire [63:0] bit_data_339,
    input wire [63:0] bit_data_340,
    input wire [63:0] bit_data_341,
    input wire [63:0] bit_data_342,
    input wire [63:0] bit_data_343,
    input wire [63:0] bit_data_344,
    input wire [63:0] bit_data_345,
    input wire [63:0] bit_data_346,
    input wire [63:0] bit_data_347,
    input wire [63:0] bit_data_348,
    input wire [63:0] bit_data_349,
    input wire [63:0] bit_data_350,
    input wire [63:0] bit_data_351,
    input wire [63:0] bit_data_352,
    input wire [63:0] bit_data_353,
    input wire [63:0] bit_data_354,
    input wire [63:0] bit_data_355,
    input wire [63:0] bit_data_356,
    input wire [63:0] bit_data_357,
    input wire [63:0] bit_data_358,
    input wire [63:0] bit_data_359,
    input wire [63:0] bit_data_360,
    input wire [63:0] bit_data_361,
    input wire [63:0] bit_data_362,
    input wire [63:0] bit_data_363,
    input wire [63:0] bit_data_364,
    input wire [63:0] bit_data_365,
    input wire [63:0] bit_data_366,
    input wire [63:0] bit_data_367,
    input wire [63:0] bit_data_368,
    input wire [63:0] bit_data_369,
    input wire [63:0] bit_data_370,
    input wire [63:0] bit_data_371,
    input wire [63:0] bit_data_372,
    input wire [63:0] bit_data_373,
    input wire [63:0] bit_data_374,
    input wire [63:0] bit_data_375,
    input wire [63:0] bit_data_376,
    input wire [63:0] bit_data_377,
    input wire [63:0] bit_data_378,
    input wire [63:0] bit_data_379,
    input wire [63:0] bit_data_380,
    input wire [63:0] bit_data_381,
    input wire [63:0] bit_data_382,
    input wire [63:0] bit_data_383,
    input wire [63:0] bit_data_384,
    input wire [63:0] bit_data_385,
    input wire [63:0] bit_data_386,
    input wire [63:0] bit_data_387,
    input wire [63:0] bit_data_388,
    input wire [63:0] bit_data_389,
    input wire [63:0] bit_data_390,
    input wire [63:0] bit_data_391,
    input wire [63:0] bit_data_392,
    input wire [63:0] bit_data_393,
    input wire [63:0] bit_data_394,
    input wire [63:0] bit_data_395,
    input wire [63:0] bit_data_396,
    input wire [63:0] bit_data_397,
    input wire [63:0] bit_data_398,
    input wire [63:0] bit_data_399,
    input wire [63:0] bit_data_400,
    input wire [63:0] bit_data_401,
    input wire [63:0] bit_data_402,
    input wire [63:0] bit_data_403,
    input wire [63:0] bit_data_404,
    input wire [63:0] bit_data_405,
    input wire [63:0] bit_data_406,
    input wire [63:0] bit_data_407,
    input wire [63:0] bit_data_408,
    input wire [63:0] bit_data_409,
    input wire [63:0] bit_data_410,
    input wire [63:0] bit_data_411,
    input wire [63:0] bit_data_412,
    input wire [63:0] bit_data_413,
    input wire [63:0] bit_data_414,
    input wire [63:0] bit_data_415,
    input wire [63:0] bit_data_416,
    input wire [63:0] bit_data_417,
    input wire [63:0] bit_data_418,
    input wire [63:0] bit_data_419,
    input wire [63:0] bit_data_420,
    input wire [63:0] bit_data_421,
    input wire [63:0] bit_data_422,
    input wire [63:0] bit_data_423,
    input wire [63:0] bit_data_424,
    input wire [63:0] bit_data_425,
    input wire [63:0] bit_data_426,
    input wire [63:0] bit_data_427,
    input wire [63:0] bit_data_428,
    input wire [63:0] bit_data_429,
    input wire [63:0] bit_data_430,
    input wire [63:0] bit_data_431,
    input wire [63:0] bit_data_432,
    input wire [63:0] bit_data_433,
    input wire [63:0] bit_data_434,
    input wire [63:0] bit_data_435,
    input wire [63:0] bit_data_436,
    input wire [63:0] bit_data_437,
    input wire [63:0] bit_data_438,
    input wire [63:0] bit_data_439,
    input wire [63:0] bit_data_440,
    input wire [63:0] bit_data_441,
    input wire [63:0] bit_data_442,
    input wire [63:0] bit_data_443,
    input wire [63:0] bit_data_444,
    input wire [63:0] bit_data_445,
    input wire [63:0] bit_data_446,
    input wire [63:0] bit_data_447,
    input wire [63:0] bit_data_448,
    input wire [63:0] bit_data_449,
    input wire [63:0] bit_data_450,
    input wire [63:0] bit_data_451,
    input wire [63:0] bit_data_452,
    input wire [63:0] bit_data_453,
    input wire [63:0] bit_data_454,
    input wire [63:0] bit_data_455,
    input wire [63:0] bit_data_456,
    input wire [63:0] bit_data_457,
    input wire [63:0] bit_data_458,
    input wire [63:0] bit_data_459,
    input wire [63:0] bit_data_460,
    input wire [63:0] bit_data_461,
    input wire [63:0] bit_data_462,
    input wire [63:0] bit_data_463,
    input wire [63:0] bit_data_464,
    input wire [63:0] bit_data_465,
    input wire [63:0] bit_data_466,
    input wire [63:0] bit_data_467,
    input wire [63:0] bit_data_468,
    input wire [63:0] bit_data_469,
    input wire [63:0] bit_data_470,
    input wire [63:0] bit_data_471,
    input wire [63:0] bit_data_472,
    input wire [63:0] bit_data_473,
    input wire [63:0] bit_data_474,
    input wire [63:0] bit_data_475,
    input wire [63:0] bit_data_476,
    input wire [63:0] bit_data_477,
    input wire [63:0] bit_data_478,
    input wire [63:0] bit_data_479,
    input wire [63:0] bit_data_480,
    input wire [63:0] bit_data_481,
    input wire [63:0] bit_data_482,
    input wire [63:0] bit_data_483,
    input wire [63:0] bit_data_484,
    input wire [63:0] bit_data_485,
    input wire [63:0] bit_data_486,
    input wire [63:0] bit_data_487,
    input wire [63:0] bit_data_488,
    input wire [63:0] bit_data_489,
    input wire [63:0] bit_data_490,
    input wire [63:0] bit_data_491,
    input wire [63:0] bit_data_492,
    input wire [63:0] bit_data_493,
    input wire [63:0] bit_data_494,
    input wire [63:0] bit_data_495,
    input wire [63:0] bit_data_496,
    input wire [63:0] bit_data_497,
    input wire [63:0] bit_data_498,
    input wire [63:0] bit_data_499,
    input wire [63:0] bit_data_500,
    input wire [63:0] bit_data_501,
    input wire [63:0] bit_data_502,
    input wire [63:0] bit_data_503,
    input wire [63:0] bit_data_504,
    input wire [63:0] bit_data_505,
    input wire [63:0] bit_data_506,
    input wire [63:0] bit_data_507,
    input wire [63:0] bit_data_508,
    input wire [63:0] bit_data_509,
    input wire [63:0] bit_data_510,
    input wire [63:0] bit_data_511,
    input wire [63:0] bit_data_512,
    input wire [63:0] bit_data_513,
    input wire [63:0] bit_data_514,
    input wire [63:0] bit_data_515,
    input wire [63:0] bit_data_516,
    input wire [63:0] bit_data_517,
    input wire [63:0] bit_data_518,
    input wire [63:0] bit_data_519,
    input wire [63:0] bit_data_520,
    input wire [63:0] bit_data_521,
    input wire [63:0] bit_data_522,
    input wire [63:0] bit_data_523,
    input wire [63:0] bit_data_524,
    input wire [63:0] bit_data_525,
    input wire [63:0] bit_data_526,
    input wire [63:0] bit_data_527,
    input wire [63:0] bit_data_528,
    input wire [63:0] bit_data_529,
    input wire [63:0] bit_data_530,
    input wire [63:0] bit_data_531,
    input wire [63:0] bit_data_532,
    input wire [63:0] bit_data_533,

        output reg [63:0] data_decode,
        output reg        data_en
    );

    // * 输出总线只需  个周期即可输出完毕
    // * 而输入总线也需要 24 个周期输出完毕，而且先计算 CFU，不会立即更新 VFU
    // * 所以没必要写入 reg 后再


    reg  [ 9:0] cnt;
    reg         flag_en;
    wire [63:0] bit_data[QC_LDPC_COL_COUNT-1:0];

    assign bit_data[0]  = bit_data_1;
    assign bit_data[1]  = bit_data_2;
    assign bit_data[2]  = bit_data_3;
    assign bit_data[3]  = bit_data_4;
    assign bit_data[4]  = bit_data_5;
    assign bit_data[5]  = bit_data_6;
    assign bit_data[6]  = bit_data_7;
    assign bit_data[7]  = bit_data_8;
    assign bit_data[8]  = bit_data_9;
    assign bit_data[9]  = bit_data_10;
    assign bit_data[10] = bit_data_11;
    assign bit_data[11] = bit_data_12;
    assign bit_data[12] = bit_data_13;
    assign bit_data[13] = bit_data_14;
    assign bit_data[14] = bit_data_15;
    assign bit_data[15] = bit_data_16;
    assign bit_data[16] = bit_data_17;
    assign bit_data[17] = bit_data_18;
    assign bit_data[18] = bit_data_19;
    assign bit_data[19] = bit_data_20;
    assign bit_data[20] = bit_data_21;
    assign bit_data[21] = bit_data_22;
    assign bit_data[22] = bit_data_23;
    assign bit_data[23] = bit_data_24;
    assign bit_data[24] = bit_data_25;
    assign bit_data[25] = bit_data_26;
    assign bit_data[26] = bit_data_27;
    assign bit_data[27] = bit_data_28;
    assign bit_data[28] = bit_data_29;
    assign bit_data[29] = bit_data_30;
    assign bit_data[30] = bit_data_31;
    assign bit_data[31] = bit_data_32;
    assign bit_data[32] = bit_data_33;
    assign bit_data[33] = bit_data_34;
    assign bit_data[34] = bit_data_35;
    assign bit_data[35] = bit_data_36;
    assign bit_data[36] = bit_data_37;
    assign bit_data[37] = bit_data_38;
    assign bit_data[38] = bit_data_39;
    assign bit_data[39] = bit_data_40;
    assign bit_data[40] = bit_data_41;
    assign bit_data[41] = bit_data_42;
    assign bit_data[42] = bit_data_43;
    assign bit_data[43] = bit_data_44;
    assign bit_data[44] = bit_data_45;
    assign bit_data[45] = bit_data_46;
    assign bit_data[46] = bit_data_47;
    assign bit_data[47] = bit_data_48;
    assign bit_data[48] = bit_data_49;
    assign bit_data[49] = bit_data_50;
    assign bit_data[50] = bit_data_51;
    assign bit_data[51] = bit_data_52;
    assign bit_data[52] = bit_data_53;
    assign bit_data[53] = bit_data_54;
    assign bit_data[54] = bit_data_55;
    assign bit_data[55] = bit_data_56;
    assign bit_data[56] = bit_data_57;
    assign bit_data[57] = bit_data_58;
    assign bit_data[58] = bit_data_59;
    assign bit_data[59] = bit_data_60;
    assign bit_data[60] = bit_data_61;
    assign bit_data[61] = bit_data_62;
    assign bit_data[62] = bit_data_63;
    assign bit_data[63] = bit_data_64;
    assign bit_data[64] = bit_data_65;
    assign bit_data[65] = bit_data_66;
    assign bit_data[66] = bit_data_67;
    assign bit_data[67] = bit_data_68;
    assign bit_data[68] = bit_data_69;
    assign bit_data[69] = bit_data_70;
    assign bit_data[70] = bit_data_71;
    assign bit_data[71] = bit_data_72;
    assign bit_data[72] = bit_data_73;
    assign bit_data[73] = bit_data_74;
    assign bit_data[74] = bit_data_75;
    assign bit_data[75] = bit_data_76;
    assign bit_data[76] = bit_data_77;
    assign bit_data[77] = bit_data_78;
    assign bit_data[78] = bit_data_79;
    assign bit_data[79] = bit_data_80;
    assign bit_data[80] = bit_data_81;
    assign bit_data[81] = bit_data_82;
    assign bit_data[82] = bit_data_83;
    assign bit_data[83] = bit_data_84;
    assign bit_data[84] = bit_data_85;
    assign bit_data[85] = bit_data_86;
    assign bit_data[86] = bit_data_87;
    assign bit_data[87] = bit_data_88;
    assign bit_data[88] = bit_data_89;
    assign bit_data[89] = bit_data_90;
    assign bit_data[90] = bit_data_91;
    assign bit_data[91] = bit_data_92;
    assign bit_data[92] = bit_data_93;
    assign bit_data[93] = bit_data_94;
    assign bit_data[94] = bit_data_95;
    assign bit_data[95] = bit_data_96;
    assign bit_data[96] = bit_data_97;
    assign bit_data[97] = bit_data_98;
    assign bit_data[98] = bit_data_99;
    assign bit_data[99] = bit_data_100;
    assign bit_data[100] = bit_data_101;
    assign bit_data[101] = bit_data_102;
    assign bit_data[102] = bit_data_103;
    assign bit_data[103] = bit_data_104;
    assign bit_data[104] = bit_data_105;
    assign bit_data[105] = bit_data_106;
    assign bit_data[106] = bit_data_107;
    assign bit_data[107] = bit_data_108;
    assign bit_data[108] = bit_data_109;
    assign bit_data[109] = bit_data_110;
    assign bit_data[110] = bit_data_111;
    assign bit_data[111] = bit_data_112;
    assign bit_data[112] = bit_data_113;
    assign bit_data[113] = bit_data_114;
    assign bit_data[114] = bit_data_115;
    assign bit_data[115] = bit_data_116;
    assign bit_data[116] = bit_data_117;
    assign bit_data[117] = bit_data_118;
    assign bit_data[118] = bit_data_119;
    assign bit_data[119] = bit_data_120;
    assign bit_data[120] = bit_data_121;
    assign bit_data[121] = bit_data_122;
    assign bit_data[122] = bit_data_123;
    assign bit_data[123] = bit_data_124;
    assign bit_data[124] = bit_data_125;
    assign bit_data[125] = bit_data_126;
    assign bit_data[126] = bit_data_127;
    assign bit_data[127] = bit_data_128;
    assign bit_data[128] = bit_data_129;
    assign bit_data[129] = bit_data_130;
    assign bit_data[130] = bit_data_131;
    assign bit_data[131] = bit_data_132;
    assign bit_data[132] = bit_data_133;
    assign bit_data[133] = bit_data_134;
    assign bit_data[134] = bit_data_135;
    assign bit_data[135] = bit_data_136;
    assign bit_data[136] = bit_data_137;
    assign bit_data[137] = bit_data_138;
    assign bit_data[138] = bit_data_139;
    assign bit_data[139] = bit_data_140;
    assign bit_data[140] = bit_data_141;
    assign bit_data[141] = bit_data_142;
    assign bit_data[142] = bit_data_143;
    assign bit_data[143] = bit_data_144;
    assign bit_data[144] = bit_data_145;
    assign bit_data[145] = bit_data_146;
    assign bit_data[146] = bit_data_147;
    assign bit_data[147] = bit_data_148;
    assign bit_data[148] = bit_data_149;
    assign bit_data[149] = bit_data_150;
    assign bit_data[150] = bit_data_151;
    assign bit_data[151] = bit_data_152;
    assign bit_data[152] = bit_data_153;
    assign bit_data[153] = bit_data_154;
    assign bit_data[154] = bit_data_155;
    assign bit_data[155] = bit_data_156;
    assign bit_data[156] = bit_data_157;
    assign bit_data[157] = bit_data_158;
    assign bit_data[158] = bit_data_159;
    assign bit_data[159] = bit_data_160;
    assign bit_data[160] = bit_data_161;
    assign bit_data[161] = bit_data_162;
    assign bit_data[162] = bit_data_163;
    assign bit_data[163] = bit_data_164;
    assign bit_data[164] = bit_data_165;
    assign bit_data[165] = bit_data_166;
    assign bit_data[166] = bit_data_167;
    assign bit_data[167] = bit_data_168;
    assign bit_data[168] = bit_data_169;
    assign bit_data[169] = bit_data_170;
    assign bit_data[170] = bit_data_171;
    assign bit_data[171] = bit_data_172;
    assign bit_data[172] = bit_data_173;
    assign bit_data[173] = bit_data_174;
    assign bit_data[174] = bit_data_175;
    assign bit_data[175] = bit_data_176;
    assign bit_data[176] = bit_data_177;
    assign bit_data[177] = bit_data_178;
    assign bit_data[178] = bit_data_179;
    assign bit_data[179] = bit_data_180;
    assign bit_data[180] = bit_data_181;
    assign bit_data[181] = bit_data_182;
    assign bit_data[182] = bit_data_183;
    assign bit_data[183] = bit_data_184;
    assign bit_data[184] = bit_data_185;
    assign bit_data[185] = bit_data_186;
    assign bit_data[186] = bit_data_187;
    assign bit_data[187] = bit_data_188;
    assign bit_data[188] = bit_data_189;
    assign bit_data[189] = bit_data_190;
    assign bit_data[190] = bit_data_191;
    assign bit_data[191] = bit_data_192;
    assign bit_data[192] = bit_data_193;
    assign bit_data[193] = bit_data_194;
    assign bit_data[194] = bit_data_195;
    assign bit_data[195] = bit_data_196;
    assign bit_data[196] = bit_data_197;
    assign bit_data[197] = bit_data_198;
    assign bit_data[198] = bit_data_199;
    assign bit_data[199] = bit_data_200;
    assign bit_data[200] = bit_data_201;
    assign bit_data[201] = bit_data_202;
    assign bit_data[202] = bit_data_203;
    assign bit_data[203] = bit_data_204;
    assign bit_data[204] = bit_data_205;
    assign bit_data[205] = bit_data_206;
    assign bit_data[206] = bit_data_207;
    assign bit_data[207] = bit_data_208;
    assign bit_data[208] = bit_data_209;
    assign bit_data[209] = bit_data_210;
    assign bit_data[210] = bit_data_211;
    assign bit_data[211] = bit_data_212;
    assign bit_data[212] = bit_data_213;
    assign bit_data[213] = bit_data_214;
    assign bit_data[214] = bit_data_215;
    assign bit_data[215] = bit_data_216;
    assign bit_data[216] = bit_data_217;
    assign bit_data[217] = bit_data_218;
    assign bit_data[218] = bit_data_219;
    assign bit_data[219] = bit_data_220;
    assign bit_data[220] = bit_data_221;
    assign bit_data[221] = bit_data_222;
    assign bit_data[222] = bit_data_223;
    assign bit_data[223] = bit_data_224;
    assign bit_data[224] = bit_data_225;
    assign bit_data[225] = bit_data_226;
    assign bit_data[226] = bit_data_227;
    assign bit_data[227] = bit_data_228;
    assign bit_data[228] = bit_data_229;
    assign bit_data[229] = bit_data_230;
    assign bit_data[230] = bit_data_231;
    assign bit_data[231] = bit_data_232;
    assign bit_data[232] = bit_data_233;
    assign bit_data[233] = bit_data_234;
    assign bit_data[234] = bit_data_235;
    assign bit_data[235] = bit_data_236;
    assign bit_data[236] = bit_data_237;
    assign bit_data[237] = bit_data_238;
    assign bit_data[238] = bit_data_239;
    assign bit_data[239] = bit_data_240;
    assign bit_data[240] = bit_data_241;
    assign bit_data[241] = bit_data_242;
    assign bit_data[242] = bit_data_243;
    assign bit_data[243] = bit_data_244;
    assign bit_data[244] = bit_data_245;
    assign bit_data[245] = bit_data_246;
    assign bit_data[246] = bit_data_247;
    assign bit_data[247] = bit_data_248;
    assign bit_data[248] = bit_data_249;
    assign bit_data[249] = bit_data_250;
    assign bit_data[250] = bit_data_251;
    assign bit_data[251] = bit_data_252;
    assign bit_data[252] = bit_data_253;
    assign bit_data[253] = bit_data_254;
    assign bit_data[254] = bit_data_255;
    assign bit_data[255] = bit_data_256;
    assign bit_data[256] = bit_data_257;
    assign bit_data[257] = bit_data_258;
    assign bit_data[258] = bit_data_259;
    assign bit_data[259] = bit_data_260;
    assign bit_data[260] = bit_data_261;
    assign bit_data[261] = bit_data_262;
    assign bit_data[262] = bit_data_263;
    assign bit_data[263] = bit_data_264;
    assign bit_data[264] = bit_data_265;
    assign bit_data[265] = bit_data_266;
    assign bit_data[266] = bit_data_267;
    assign bit_data[267] = bit_data_268;
    assign bit_data[268] = bit_data_269;
    assign bit_data[269] = bit_data_270;
    assign bit_data[270] = bit_data_271;
    assign bit_data[271] = bit_data_272;
    assign bit_data[272] = bit_data_273;
    assign bit_data[273] = bit_data_274;
    assign bit_data[274] = bit_data_275;
    assign bit_data[275] = bit_data_276;
    assign bit_data[276] = bit_data_277;
    assign bit_data[277] = bit_data_278;
    assign bit_data[278] = bit_data_279;
    assign bit_data[279] = bit_data_280;
    assign bit_data[280] = bit_data_281;
    assign bit_data[281] = bit_data_282;
    assign bit_data[282] = bit_data_283;
    assign bit_data[283] = bit_data_284;
    assign bit_data[284] = bit_data_285;
    assign bit_data[285] = bit_data_286;
    assign bit_data[286] = bit_data_287;
    assign bit_data[287] = bit_data_288;
    assign bit_data[288] = bit_data_289;
    assign bit_data[289] = bit_data_290;
    assign bit_data[290] = bit_data_291;
    assign bit_data[291] = bit_data_292;
    assign bit_data[292] = bit_data_293;
    assign bit_data[293] = bit_data_294;
    assign bit_data[294] = bit_data_295;
    assign bit_data[295] = bit_data_296;
    assign bit_data[296] = bit_data_297;
    assign bit_data[297] = bit_data_298;
    assign bit_data[298] = bit_data_299;
    assign bit_data[299] = bit_data_300;
    assign bit_data[300] = bit_data_301;
    assign bit_data[301] = bit_data_302;
    assign bit_data[302] = bit_data_303;
    assign bit_data[303] = bit_data_304;
    assign bit_data[304] = bit_data_305;
    assign bit_data[305] = bit_data_306;
    assign bit_data[306] = bit_data_307;
    assign bit_data[307] = bit_data_308;
    assign bit_data[308] = bit_data_309;
    assign bit_data[309] = bit_data_310;
    assign bit_data[310] = bit_data_311;
    assign bit_data[311] = bit_data_312;
    assign bit_data[312] = bit_data_313;
    assign bit_data[313] = bit_data_314;
    assign bit_data[314] = bit_data_315;
    assign bit_data[315] = bit_data_316;
    assign bit_data[316] = bit_data_317;
    assign bit_data[317] = bit_data_318;
    assign bit_data[318] = bit_data_319;
    assign bit_data[319] = bit_data_320;
    assign bit_data[320] = bit_data_321;
    assign bit_data[321] = bit_data_322;
    assign bit_data[322] = bit_data_323;
    assign bit_data[323] = bit_data_324;
    assign bit_data[324] = bit_data_325;
    assign bit_data[325] = bit_data_326;
    assign bit_data[326] = bit_data_327;
    assign bit_data[327] = bit_data_328;
    assign bit_data[328] = bit_data_329;
    assign bit_data[329] = bit_data_330;
    assign bit_data[330] = bit_data_331;
    assign bit_data[331] = bit_data_332;
    assign bit_data[332] = bit_data_333;
    assign bit_data[333] = bit_data_334;
    assign bit_data[334] = bit_data_335;
    assign bit_data[335] = bit_data_336;
    assign bit_data[336] = bit_data_337;
    assign bit_data[337] = bit_data_338;
    assign bit_data[338] = bit_data_339;
    assign bit_data[339] = bit_data_340;
    assign bit_data[340] = bit_data_341;
    assign bit_data[341] = bit_data_342;
    assign bit_data[342] = bit_data_343;
    assign bit_data[343] = bit_data_344;
    assign bit_data[344] = bit_data_345;
    assign bit_data[345] = bit_data_346;
    assign bit_data[346] = bit_data_347;
    assign bit_data[347] = bit_data_348;
    assign bit_data[348] = bit_data_349;
    assign bit_data[349] = bit_data_350;
    assign bit_data[350] = bit_data_351;
    assign bit_data[351] = bit_data_352;
    assign bit_data[352] = bit_data_353;
    assign bit_data[353] = bit_data_354;
    assign bit_data[354] = bit_data_355;
    assign bit_data[355] = bit_data_356;
    assign bit_data[356] = bit_data_357;
    assign bit_data[357] = bit_data_358;
    assign bit_data[358] = bit_data_359;
    assign bit_data[359] = bit_data_360;
    assign bit_data[360] = bit_data_361;
    assign bit_data[361] = bit_data_362;
    assign bit_data[362] = bit_data_363;
    assign bit_data[363] = bit_data_364;
    assign bit_data[364] = bit_data_365;
    assign bit_data[365] = bit_data_366;
    assign bit_data[366] = bit_data_367;
    assign bit_data[367] = bit_data_368;
    assign bit_data[368] = bit_data_369;
    assign bit_data[369] = bit_data_370;
    assign bit_data[370] = bit_data_371;
    assign bit_data[371] = bit_data_372;
    assign bit_data[372] = bit_data_373;
    assign bit_data[373] = bit_data_374;
    assign bit_data[374] = bit_data_375;
    assign bit_data[375] = bit_data_376;
    assign bit_data[376] = bit_data_377;
    assign bit_data[377] = bit_data_378;
    assign bit_data[378] = bit_data_379;
    assign bit_data[379] = bit_data_380;
    assign bit_data[380] = bit_data_381;
    assign bit_data[381] = bit_data_382;
    assign bit_data[382] = bit_data_383;
    assign bit_data[383] = bit_data_384;
    assign bit_data[384] = bit_data_385;
    assign bit_data[385] = bit_data_386;
    assign bit_data[386] = bit_data_387;
    assign bit_data[387] = bit_data_388;
    assign bit_data[388] = bit_data_389;
    assign bit_data[389] = bit_data_390;
    assign bit_data[390] = bit_data_391;
    assign bit_data[391] = bit_data_392;
    assign bit_data[392] = bit_data_393;
    assign bit_data[393] = bit_data_394;
    assign bit_data[394] = bit_data_395;
    assign bit_data[395] = bit_data_396;
    assign bit_data[396] = bit_data_397;
    assign bit_data[397] = bit_data_398;
    assign bit_data[398] = bit_data_399;
    assign bit_data[399] = bit_data_400;
    assign bit_data[400] = bit_data_401;
    assign bit_data[401] = bit_data_402;
    assign bit_data[402] = bit_data_403;
    assign bit_data[403] = bit_data_404;
    assign bit_data[404] = bit_data_405;
    assign bit_data[405] = bit_data_406;
    assign bit_data[406] = bit_data_407;
    assign bit_data[407] = bit_data_408;
    assign bit_data[408] = bit_data_409;
    assign bit_data[409] = bit_data_410;
    assign bit_data[410] = bit_data_411;
    assign bit_data[411] = bit_data_412;
    assign bit_data[412] = bit_data_413;
    assign bit_data[413] = bit_data_414;
    assign bit_data[414] = bit_data_415;
    assign bit_data[415] = bit_data_416;
    assign bit_data[416] = bit_data_417;
    assign bit_data[417] = bit_data_418;
    assign bit_data[418] = bit_data_419;
    assign bit_data[419] = bit_data_420;
    assign bit_data[420] = bit_data_421;
    assign bit_data[421] = bit_data_422;
    assign bit_data[422] = bit_data_423;
    assign bit_data[423] = bit_data_424;
    assign bit_data[424] = bit_data_425;
    assign bit_data[425] = bit_data_426;
    assign bit_data[426] = bit_data_427;
    assign bit_data[427] = bit_data_428;
    assign bit_data[428] = bit_data_429;
    assign bit_data[429] = bit_data_430;
    assign bit_data[430] = bit_data_431;
    assign bit_data[431] = bit_data_432;
    assign bit_data[432] = bit_data_433;
    assign bit_data[433] = bit_data_434;
    assign bit_data[434] = bit_data_435;
    assign bit_data[435] = bit_data_436;
    assign bit_data[436] = bit_data_437;
    assign bit_data[437] = bit_data_438;
    assign bit_data[438] = bit_data_439;
    assign bit_data[439] = bit_data_440;
    assign bit_data[440] = bit_data_441;
    assign bit_data[441] = bit_data_442;
    assign bit_data[442] = bit_data_443;
    assign bit_data[443] = bit_data_444;
    assign bit_data[444] = bit_data_445;
    assign bit_data[445] = bit_data_446;
    assign bit_data[446] = bit_data_447;
    assign bit_data[447] = bit_data_448;
    assign bit_data[448] = bit_data_449;
    assign bit_data[449] = bit_data_450;
    assign bit_data[450] = bit_data_451;
    assign bit_data[451] = bit_data_452;
    assign bit_data[452] = bit_data_453;
    assign bit_data[453] = bit_data_454;
    assign bit_data[454] = bit_data_455;
    assign bit_data[455] = bit_data_456;
    assign bit_data[456] = bit_data_457;
    assign bit_data[457] = bit_data_458;
    assign bit_data[458] = bit_data_459;
    assign bit_data[459] = bit_data_460;
    assign bit_data[460] = bit_data_461;
    assign bit_data[461] = bit_data_462;
    assign bit_data[462] = bit_data_463;
    assign bit_data[463] = bit_data_464;
    assign bit_data[464] = bit_data_465;
    assign bit_data[465] = bit_data_466;
    assign bit_data[466] = bit_data_467;
    assign bit_data[467] = bit_data_468;
    assign bit_data[468] = bit_data_469;
    assign bit_data[469] = bit_data_470;
    assign bit_data[470] = bit_data_471;
    assign bit_data[471] = bit_data_472;
    assign bit_data[472] = bit_data_473;
    assign bit_data[473] = bit_data_474;
    assign bit_data[474] = bit_data_475;
    assign bit_data[475] = bit_data_476;
    assign bit_data[476] = bit_data_477;
    assign bit_data[477] = bit_data_478;
    assign bit_data[478] = bit_data_479;
    assign bit_data[479] = bit_data_480;
    assign bit_data[480] = bit_data_481;
    assign bit_data[481] = bit_data_482;
    assign bit_data[482] = bit_data_483;
    assign bit_data[483] = bit_data_484;
    assign bit_data[484] = bit_data_485;
    assign bit_data[485] = bit_data_486;
    assign bit_data[486] = bit_data_487;
    assign bit_data[487] = bit_data_488;
    assign bit_data[488] = bit_data_489;
    assign bit_data[489] = bit_data_490;
    assign bit_data[490] = bit_data_491;
    assign bit_data[491] = bit_data_492;
    assign bit_data[492] = bit_data_493;
    assign bit_data[493] = bit_data_494;
    assign bit_data[494] = bit_data_495;
    assign bit_data[495] = bit_data_496;
    assign bit_data[496] = bit_data_497;
    assign bit_data[497] = bit_data_498;
    assign bit_data[498] = bit_data_499;
    assign bit_data[499] = bit_data_500;
    assign bit_data[500] = bit_data_501;
    assign bit_data[501] = bit_data_502;
    assign bit_data[502] = bit_data_503;
    assign bit_data[503] = bit_data_504;
    assign bit_data[504] = bit_data_505;
    assign bit_data[505] = bit_data_506;
    assign bit_data[506] = bit_data_507;
    assign bit_data[507] = bit_data_508;
    assign bit_data[508] = bit_data_509;
    assign bit_data[509] = bit_data_510;
    assign bit_data[510] = bit_data_511;
    assign bit_data[511] = bit_data_512;
    assign bit_data[512] = bit_data_513;
    assign bit_data[513] = bit_data_514;
    assign bit_data[514] = bit_data_515;
    assign bit_data[515] = bit_data_516;
    assign bit_data[516] = bit_data_517;
    assign bit_data[517] = bit_data_518;
    assign bit_data[518] = bit_data_519;
    assign bit_data[519] = bit_data_520;
    assign bit_data[520] = bit_data_521;
    assign bit_data[521] = bit_data_522;
    assign bit_data[522] = bit_data_523;
    assign bit_data[523] = bit_data_524;
    assign bit_data[524] = bit_data_525;
    assign bit_data[525] = bit_data_526;
    assign bit_data[526] = bit_data_527;
    assign bit_data[527] = bit_data_528;
    assign bit_data[528] = bit_data_529;
    assign bit_data[529] = bit_data_530;
    assign bit_data[530] = bit_data_531;
    assign bit_data[531] = bit_data_532;
    assign bit_data[532] = bit_data_533;




    // 输出地址计数器
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            cnt <= 10'd0;
        else if (cnt == QC_LDPC_COL_COUNT - 1)
            cnt <= 10'd0;
        else if (flag_en == 1'b1)
            cnt <= cnt + 1'b1;
        else
            cnt <= cnt;

    // 将一个周期的 en 信号扩展为 127 个周期
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            flag_en <= 1'b0;
        else if (cnt == QC_LDPC_COL_COUNT - 1)
            flag_en <= 1'b0;
        else if (flag_serial == 1'b1)
            flag_en <= 1'b1;
        else
            flag_en <= flag_en;

    // 给 flag_en 打一拍以实现控制与数据的同步
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            data_en <= 1'b0;
        else
            data_en <= flag_en;

    // 硬判决数据结果输出，但是因为连线的时候没有从 0 开始，故进行 cnt+1'b1
    always @(posedge sys_clk or negedge sys_rst_n)
        if (sys_rst_n == 1'b0)
            data_decode <= 64'd0;
        else if (flag_en == 1'b1)
            data_decode <= bit_data[cnt];
        else
            data_decode <= 64'dz;
endmodule
